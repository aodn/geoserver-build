netcdf file-91.nc {
  dimensions:
    DEPTH = 21;
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073, 23178.750011574073}
TEMP =
  {27.0045, 27.0286, 27.0308, 27.0324, 27.0317, 27.0298, 27.0325, 27.0356, 27.0365, 27.0368, 27.0365, 27.0359, 27.0359, 27.0365, 27.0351, 27.0325, 27.0311, 27.0304, 27.0321, 27.0344, 27.0346}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872}
}
