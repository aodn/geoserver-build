netcdf file-82.nc {
  dimensions:
    DEPTH = 20;
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406, 23178.419907407406}
TEMP =
  {26.9885, 26.9894, 26.9902, 26.9928, 26.9951, 26.997, 26.9998, 26.9996, 26.9986, 26.9999, 27.0, 27.0013, 27.0023, 27.0023, 27.002, 27.0027, 27.003, 27.0026, 27.0027, 27.0037}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.908, 15.903, 16.897, 17.89, 18.884, 19.878}
}
