netcdf file-11.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (48 currently)
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875, 22509.1221875}
TEMP =
  {16.3794, 16.3609, 16.3543, 16.3511, 16.3493, 16.3488, 16.3464, 16.3447, 16.3427, 16.3424, 16.3425, 16.341, 16.3386, 16.3374, 16.3364, 16.3326, 16.3294, 16.3222, 16.3078, 16.3019, 16.2912, 16.2775, 16.2667, 16.2613, 16.2558, 16.2485, 16.2456, 16.244, 16.2427, 16.2417, 16.2415, 16.2414, 16.2412, 16.2404, 16.2365, 16.234, 16.2334, 16.2333, 16.2335, 16.2338, 16.2341, 16.2342, 16.2348, 16.2359, 16.2363, 16.236, 16.2355, 16.2354}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0}
}
