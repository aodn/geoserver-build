netcdf file-149.nc {
  dimensions:
    DEPTH = 25;
  variables:
    float LATITUDE(DEPTH=25);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=25);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=25);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=25);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=25);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=25);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593, 21898.071030092593}
TEMP =
  {27.4866, 27.5359, 27.5381, 27.5288, 27.5146, 27.5149, 27.5127, 27.5112, 27.5094, 27.5064, 27.5046, 27.5033, 27.503, 27.5016, 27.5001, 27.4994, 27.4988, 27.4984, 27.4979, 27.497, 27.4967, 27.497, 27.4971, 27.4975, 27.4977}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.902, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847}
}
