netcdf file-37.nc {
  dimensions:
    DEPTH = 43;
  variables:
    float LATITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=43);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=43);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741, 22304.07115740741}
TEMP =
  {22.401, 22.3991, 22.3951, 22.3947, 22.3941, 22.394, 22.3945, 22.3937, 22.3961, 22.403, 22.4095, 22.4108, 22.3993, 22.3848, 22.3616, 22.2736, 22.1995, 22.126, 22.0898, 22.0685, 22.0593, 22.0494, 22.049, 22.0478, 22.0454, 22.0404, 22.0245, 21.9949, 21.9614, 21.9397, 21.9156, 21.8859, 21.8283, 21.7515, 21.6293, 21.4995, 21.473, 21.4439, 21.4101, 21.3794, 21.3703, 21.3732, 21.3722}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
