netcdf file-118.nc {
  dimensions:
    DEPTH = 19;
  variables:
    float LATITUDE(DEPTH=19);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=19);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=19);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=19);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=19);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=19);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98, 22987.98}
TEMP =
  {31.899, 31.8963, 31.8957, 31.8952, 31.8948, 31.894, 31.8893, 31.888, 31.8886, 31.8852, 31.8831, 31.8813, 31.8813, 31.8814, 31.8816, 31.8822, 31.8826, 31.882, 31.8809}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884}
}
