netcdf file-38.nc {
  dimensions:
    DEPTH = 45;
  variables:
    float LATITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=45);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=45);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964, 22334.080775462964}
TEMP =
  {24.6132, 24.6237, 24.5864, 24.5532, 24.5479, 24.5567, 24.5401, 24.5201, 24.5135, 24.5066, 24.5017, 24.5007, 24.5042, 24.4967, 24.4905, 24.4839, 24.453, 24.3693, 24.3004, 24.255, 24.2037, 24.1896, 24.1905, 24.1853, 24.1835, 24.184, 24.1861, 24.1905, 24.1892, 24.1898, 24.1862, 24.1834, 24.1854, 24.1834, 24.1803, 24.1794, 24.1763, 24.176, 24.1757, 24.1749, 24.1736, 24.1724, 24.1723, 24.1708, 24.1703}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
