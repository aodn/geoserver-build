netcdf file-164.nc {
  dimensions:
    DEPTH = 11;
  variables:
    float LATITUDE(DEPTH=11);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=11);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=11);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=11);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=11);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=11);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963, 22502.04712962963}
TEMP =
  {21.7919, 21.8274, 21.8575, 21.8776, 21.8866, 21.8905, 21.8919, 21.8928, 21.8941, 21.8954, 21.8976}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.854, 24.847, 25.841, 26.835}
}
