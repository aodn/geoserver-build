netcdf file-33.nc {
  dimensions:
    DEPTH = 40;
  variables:
    float LATITUDE(DEPTH=40);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=40);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=40);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=40);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=40);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=40);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925, 22150.310925925925}
TEMP =
  {20.2709, 20.5149, 20.525, 20.5252, 20.5245, 20.5226, 20.5162, 20.493, 20.4401, 20.3458, 20.2456, 20.1833, 20.1318, 20.0391, 19.9166, 19.8813, 19.856, 19.8374, 19.8436, 19.8647, 19.8812, 19.8178, 19.7089, 19.5869, 19.0969, 18.3656, 18.0927, 18.0431, 18.0322, 18.0282, 18.0269, 18.0256, 18.0239, 18.0232, 18.0231, 18.0237, 18.0223, 18.018, 18.015, 18.011}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0}
}
