netcdf file-48.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (46 currently)
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963, 22733.07994212963}
TEMP =
  {23.0598, 22.9978, 22.9754, 22.972, 22.971, 22.9695, 22.9712, 22.9707, 22.9726, 22.9706, 22.9699, 22.9751, 22.976, 22.9708, 22.9632, 22.935, 22.9226, 22.9256, 22.9202, 22.9132, 22.9115, 22.9109, 22.9107, 22.9088, 22.9086, 22.9078, 22.905, 22.9048, 22.903, 22.8992, 22.8962, 22.8952, 22.8924, 22.8916, 22.892, 22.8924, 22.8932, 22.893, 22.8923, 22.8929, 22.8936, 22.8942, 22.895, 22.894, 22.8931, 22.8937}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
