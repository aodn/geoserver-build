netcdf file-18.nc {
  dimensions:
    DEPTH = 48;
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334, -33.933334}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148, 23083.07898148148}
TEMP =
  {21.1669, 21.1665, 21.1639, 21.1591, 21.1542, 21.1513, 21.1487, 21.1477, 21.1473, 21.1472, 21.1471, 21.1484, 21.1489, 21.1484, 21.1479, 21.1476, 21.1452, 21.1443, 21.1435, 21.1429, 21.1423, 21.1426, 21.1423, 21.1434, 21.1441, 21.1446, 21.1449, 21.1431, 21.1404, 21.1402, 21.1402, 21.1405, 21.1409, 21.1406, 21.1408, 21.1406, 21.1407, 21.1405, 21.139, 21.1394, 21.1388, 21.1381, 21.1384, 21.1394, 21.1398, 21.1402, 21.1406, 21.141}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
