netcdf file-72.nc {
  dimensions:
    DEPTH = 44;
  variables:
    float LATITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=44);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=44);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704, 22634.32859953704}
TEMP =
  {22.119205, 22.1171, 22.115116, 22.114353, 22.11301, 22.104582, 22.09533, 22.0788, 22.080223, 22.020737, 21.883797, 21.83421, 21.80694, 21.78281, 21.76185, 21.73695, 21.664112, 21.591919, 21.583607, 21.572641, 21.555082, 21.511316, 21.507442, 21.50516, 21.500124, 21.498865, 21.495594, 21.487854, 21.46474, 21.444939, 21.403954, 21.345856, 21.338587, 21.326258, 21.321377, 21.312305, 21.304827, 21.297138, 21.292791, 21.286957, 21.161375, 21.028404, 20.77519, 20.728493}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0}
}
