netcdf file-100.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778, 22658.93934027778}
TEMP =
  {31.4858, 31.4893, 31.4885, 31.4897, 31.4905, 31.4892, 31.486, 31.4816, 31.4786, 31.4764, 31.4741, 31.4712, 31.469, 31.467, 31.4644, 31.4593, 31.4512, 31.4463, 31.4443, 31.443, 31.4419}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.989, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.949, 9.942, 10.936, 11.931, 12.926, 13.92, 14.914, 15.908, 16.902, 17.897, 18.891, 19.885, 20.879}
}
