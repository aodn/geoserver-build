netcdf file-110.nc {
  dimensions:
    DEPTH = 22;
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037, 22987.68818287037}
TEMP =
  {31.922, 31.9209, 31.9216, 31.9219, 31.9218, 31.9219, 31.9234, 31.9253, 31.926, 31.9247, 31.918, 31.9079, 31.9045, 31.9042, 31.9048, 31.9062, 31.9067, 31.9062, 31.9057, 31.9058, 31.9064, 31.9068}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879, 21.873, 22.867}
}
