netcdf file-102.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (20 currently)
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148, 22659.02335648148}
TEMP =
  {31.4196, 31.4202, 31.427, 31.4326, 31.4361, 31.4371, 31.4365, 31.436, 31.4352, 31.4329, 31.4308, 31.4297, 31.4286, 31.428, 31.426, 31.4231, 31.4216, 31.4206, 31.4198, 31.4197}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.891, 19.885, 20.879, 21.873, 22.867}
}
