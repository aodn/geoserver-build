netcdf file-16.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (49 currently)
  variables:
    float LATITUDE(DEPTH=49);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=49);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=49);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=49);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=49);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=49);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667, -33.931667}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927, 22898.238738425927}
TEMP =
  {16.5675, 16.5738, 16.5729, 16.5736, 16.5738, 16.5729, 16.5723, 16.5657, 16.5577, 16.5525, 16.5534, 16.5501, 16.542, 16.536, 16.5314, 16.5271, 16.5246, 16.5228, 16.5182, 16.5137, 16.5056, 16.5009, 16.4986, 16.4948, 16.489, 16.4833, 16.4628, 16.4528, 16.4489, 16.4467, 16.4423, 16.4342, 16.4246, 16.4168, 16.4034, 16.3767, 16.3311, 16.2889, 16.2668, 16.2519, 16.2413, 16.2369, 16.232, 16.2226, 16.2098, 16.1945, 16.1866, 16.1787, 16.1741}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0}
}
