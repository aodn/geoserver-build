netcdf file-125.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (25 currently)
  variables:
    float LATITUDE(DEPTH=25);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=25);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=25);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=25);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=25);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=25);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667, 22906.048854166667}
TEMP =
  {23.8754, 23.8148, 23.73, 23.6601, 23.6086, 23.5869, 23.5731, 23.5584, 23.5176, 23.4671, 23.4417, 23.4273, 23.421, 23.4165, 23.4122, 23.4081, 23.4077, 23.407, 23.4065, 23.4053, 23.4054, 23.4053, 23.4056, 23.4059, 23.4051}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847}
}
