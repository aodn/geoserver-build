netcdf file-174.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (27 currently)
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854, 22873.066226851854}
TEMP =
  {21.7075, 21.6937, 21.6817, 21.685, 21.6734, 21.6661, 21.6598, 21.6487, 21.6411, 21.6365, 21.626, 21.6235, 21.625, 21.6146, 21.6132, 21.6128, 21.613, 21.6133, 21.6136, 21.6137, 21.6134, 21.6124, 21.6123, 21.6131, 21.6133, 21.616, 21.6234}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.854, 24.847, 25.841, 26.835, 27.829}
}
