netcdf file-170.nc {
  dimensions:
    DEPTH = 28;
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147, 22737.043773148147}
TEMP =
  {27.6804, 27.7069, 27.662, 27.6343, 27.6167, 27.604, 27.5949, 27.5886, 27.5838, 27.5803, 27.5777, 27.5754, 27.5733, 27.5714, 27.5701, 27.5692, 27.5686, 27.5683, 27.5682, 27.5681, 27.5683, 27.5683, 27.5684, 27.5686, 27.5688, 27.5692, 27.5698, 27.5703}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.993, 1.989, 2.982, 3.975, 4.969, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.828}
}
