netcdf file-169.nc {
  dimensions:
    DEPTH = 30;
  variables:
    float LATITUDE(DEPTH=30);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=30);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=30);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=30);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=30);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=30);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443, 22683.051319444443}
TEMP =
  {29.7665, 29.7485, 29.725, 29.6577, 29.5786, 29.5382, 29.5039, 29.4657, 29.4421, 29.4268, 29.4122, 29.3657, 29.2092, 28.9716, 28.7754, 28.6789, 28.6321, 28.6036, 28.5862, 28.5773, 28.5727, 28.5702, 28.5686, 28.5676, 28.5674, 28.5672, 28.5665, 28.5663, 28.5665, 28.5669}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829, 28.823, 29.816}
}
