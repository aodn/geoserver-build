netcdf file-17.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (47 currently)
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185, 22991.094247685185}
TEMP =
  {19.6218, 19.2023, 19.3772, 19.3742, 19.3741, 19.3719, 19.3688, 19.3659, 19.3657, 19.3708, 19.3696, 19.3631, 19.3498, 19.3498, 19.3284, 19.311, 19.2997, 19.2851, 19.2589, 19.238, 19.2305, 19.207, 19.1605, 19.1027, 19.0325, 18.9584, 18.9072, 18.8849, 18.8725, 18.8584, 18.8071, 18.7332, 18.6775, 18.6531, 18.6454, 18.6432, 18.6421, 18.6413, 18.6405, 18.64, 18.6395, 18.6391, 18.6389, 18.639, 18.6392, 18.6391, 18.6392}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
