netcdf file-94.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815, 23178.828252314815}
TEMP =
  {26.7855, 27.0982, 26.9628, 26.9633, 26.9624, 26.9615, 26.9645, 26.9706, 26.9732, 26.9735, 26.9725, 26.9719, 26.9705, 26.9692, 26.9686, 26.9698, 26.9684, 26.9637, 26.9582, 26.9554, 26.9545}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.992, 1.99, 2.982, 3.976, 4.97, 5.963, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.908, 15.902, 16.896, 17.89, 18.884, 19.878, 20.872}
}
