netcdf file-46.nc {
  dimensions:
    DEPTH = 46;
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038, 22605.316099537038}
TEMP =
  {20.9846, 20.9723, 20.9264, 20.8064, 20.6372, 20.5767, 20.555, 20.5397, 20.5245, 20.5104, 20.4935, 20.4779, 20.4595, 20.4409, 20.425, 20.4169, 20.4092, 20.4026, 20.3973, 20.3884, 20.3813, 20.3772, 20.3738, 20.3723, 20.3712, 20.3702, 20.3694, 20.3653, 20.3603, 20.3576, 20.3554, 20.3519, 20.3497, 20.347, 20.3428, 20.3405, 20.3096, 20.1393, 19.8833, 19.5524, 19.3774, 19.2037, 19.0545, 18.9933, 18.9839, 18.9819}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
