netcdf file-3.nc {
  dimensions:
    DEPTH = 46;
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875, 21723.37875}
TEMP =
  {17.5368, 17.5464, 17.5504, 17.5505, 17.5504, 17.553, 17.5555, 17.5564, 17.5567, 17.5575, 17.5589, 17.5615, 17.563, 17.5628, 17.5631, 17.5638, 17.5644, 17.5647, 17.5646, 17.5646, 17.5647, 17.5642, 17.5631, 17.5611, 17.5589, 17.5564, 17.5539, 17.5522, 17.5508, 17.5495, 17.5486, 17.5477, 17.546, 17.5429, 17.5408, 17.5396, 17.5362, 17.5316, 17.528, 17.523, 17.5189, 17.5153, 17.5083, 17.501, 17.4954, 17.4916}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
