netcdf file-131.nc {
  dimensions:
    DEPTH = 28;
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444, 23145.025381944444}
TEMP =
  {25.1338, 25.1303, 25.1236, 25.1159, 25.1118, 25.1101, 25.1094, 25.1086, 25.1077, 25.1079, 25.1109, 25.1137, 25.1269, 25.1589, 25.2031, 25.2504, 25.2828, 25.3164, 25.3486, 25.3699, 25.3807, 25.3864, 25.3891, 25.3901, 25.3904, 25.3908, 25.3916, 25.3921}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
