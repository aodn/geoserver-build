netcdf file-101.nc {
  dimensions:
    DEPTH = 23;
  variables:
    float LATITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=23);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=23);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852, 22658.98039351852}
TEMP =
  {31.3699, 31.3798, 31.3841, 31.3871, 31.3961, 31.3997, 31.4066, 31.4142, 31.4148, 31.415, 31.4161, 31.4178, 31.4188, 31.4207, 31.4201, 31.4201, 31.4216, 31.421, 31.4205, 31.4228, 31.4272, 31.4299, 31.4312}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89, 19.885, 20.879, 21.873, 22.867}
}
