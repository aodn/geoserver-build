netcdf file-127.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (28 currently)
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926, 22978.03332175926}
TEMP =
  {27.1792, 27.1716, 27.1504, 27.1194, 27.1035, 27.0963, 27.0943, 27.0931, 27.0926, 27.0921, 27.091, 27.0886, 27.0852, 27.081, 27.0771, 27.0766, 27.081, 27.0814, 27.0791, 27.0773, 27.0784, 27.0773, 27.0768, 27.0768, 27.077, 27.0773, 27.0776, 27.078}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.891, 18.885, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
