netcdf file-107.nc {
  dimensions:
    DEPTH = 20;
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111, 22659.23048611111}
TEMP =
  {31.5523, 31.554, 31.5542, 31.5541, 31.5558, 31.5543, 31.5509, 31.5476, 31.5459, 31.5445, 31.5441, 31.5435, 31.5435, 31.5436, 31.5433, 31.5434, 31.5438, 31.544, 31.5439, 31.5439}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.989, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89, 19.885}
}
