netcdf file-14.nc {
  dimensions:
    DEPTH = 50;
  variables:
    float LATITUDE(DEPTH=50);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=50);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=50);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=50);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=50);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=50);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074, 22713.07542824074}
TEMP =
  {20.8462, 20.8473, 20.845, 20.8413, 20.8403, 20.8376, 20.8372, 20.8364, 20.8359, 20.8355, 20.8339, 20.8302, 20.8298, 20.8297, 20.8294, 20.8296, 20.8288, 20.8285, 20.8276, 20.8288, 20.8307, 20.8308, 20.8294, 20.8278, 20.8264, 20.8275, 20.8307, 20.8306, 20.831, 20.8313, 20.8349, 20.8373, 20.836, 20.8343, 20.8363, 20.8342, 20.8324, 20.8328, 20.8333, 20.8342, 20.8345, 20.833, 20.8311, 20.8361, 20.8425, 20.8466, 20.8429, 20.8405, 20.8345, 20.8352}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0}
}
