netcdf file-163.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (16 currently)
  variables:
    float LATITUDE(DEPTH=16);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=16);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=16);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=16);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=16);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=16);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964, 22480.095775462964}
TEMP =
  {21.723, 21.7202, 21.7177, 21.7163, 21.7154, 21.7145, 21.7129, 21.7118, 21.7115, 21.7116, 21.7118, 21.7121, 21.7125, 21.7126, 21.7129, 21.713}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847}
}
