netcdf file-152.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (22 currently)
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778, 22017.17809027778}
TEMP =
  {27.2914, 27.3416, 27.3727, 27.389, 27.3899, 27.3905, 27.3906, 27.3904, 27.3903, 27.3903, 27.3904, 27.3906, 27.3908, 27.3907, 27.3902, 27.3918, 27.3923, 27.3929, 27.3934, 27.3943, 27.3952, 27.3972}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.891, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
