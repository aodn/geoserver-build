netcdf IMOS_ANMN-TS_20150113T230000Z_WATR20_FV01_WATR20-1407-Seabird-SBE39-600m-temp-only-100_END-20150121T032000Z_id-7737.nc {
  dimensions:
    TIME = 1035;
  variables:
    double TIME(TIME=1035);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=1035);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=1035);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=1035);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=1035);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=1035);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=1035);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=1035);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=1035);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=1035);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=1035);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=1035);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=1035);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been filled using the DEPTH median (mooring).";
  :instrument = "Seabird         SBE39 [600m] temp only";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "3949303-4125";
  :history = "2015-01-29T06:32:01Z - depthPP: Depth computed from the 2 nearest pressure sensors available, using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 100.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = 0.0703091f; // float
  :geospatial_vertical_max = 111.37032f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-21T03:20:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.965277777777, 23753.972222222223, 23753.979166666668, 23753.98611111111, 23753.993055555555, 23754.0, 23754.006944444445, 23754.01388888889, 23754.020833333332, 23754.027777777777, 23754.034722222223, 23754.041666666668, 23754.04861111111, 23754.055555555555, 23754.0625, 23754.069444444445, 23754.07638888889, 23754.083333333332, 23754.090277777777, 23754.097222222223, 23754.104166666668, 23754.11111111111, 23754.118055555555, 23754.125, 23754.131944444445, 23754.13888888889, 23754.145833333332, 23754.152777777777, 23754.159722222223, 23754.166666666668, 23754.17361111111, 23754.180555555555, 23754.1875, 23754.194444444445, 23754.20138888889, 23754.208333333332, 23754.215277777777, 23754.222222222223, 23754.229166666668, 23754.23611111111, 23754.243055555555, 23754.25, 23754.256944444445, 23754.26388888889, 23754.270833333332, 23754.277777777777, 23754.284722222223, 23754.291666666668, 23754.29861111111, 23754.305555555555, 23754.3125, 23754.319444444445, 23754.32638888889, 23754.333333333332, 23754.340277777777, 23754.347222222223, 23754.354166666668, 23754.36111111111, 23754.368055555555, 23754.375, 23754.381944444445, 23754.38888888889, 23754.395833333332, 23754.402777777777, 23754.409722222223, 23754.416666666668, 23754.42361111111, 23754.430555555555, 23754.4375, 23754.444444444445, 23754.45138888889, 23754.458333333332, 23754.465277777777, 23754.472222222223, 23754.479166666668, 23754.48611111111, 23754.493055555555, 23754.5, 23754.506944444445, 23754.51388888889, 23754.520833333332, 23754.527777777777, 23754.534722222223, 23754.541666666668, 23754.54861111111, 23754.555555555555, 23754.5625, 23754.569444444445, 23754.57638888889, 23754.583333333332, 23754.590277777777, 23754.597222222223, 23754.604166666668, 23754.61111111111, 23754.618055555555, 23754.625, 23754.631944444445, 23754.63888888889, 23754.645833333332, 23754.652777777777, 23754.659722222223, 23754.666666666668, 23754.67361111111, 23754.680555555555, 23754.6875, 23754.694444444445, 23754.70138888889, 23754.708333333332, 23754.715277777777, 23754.722222222223, 23754.729166666668, 23754.73611111111, 23754.743055555555, 23754.75, 23754.756944444445, 23754.76388888889, 23754.770833333332, 23754.777777777777, 23754.784722222223, 23754.791666666668, 23754.79861111111, 23754.805555555555, 23754.8125, 23754.819444444445, 23754.82638888889, 23754.833333333332, 23754.840277777777, 23754.847222222223, 23754.854166666668, 23754.86111111111, 23754.868055555555, 23754.875, 23754.881944444445, 23754.88888888889, 23754.895833333332, 23754.902777777777, 23754.909722222223, 23754.916666666668, 23754.92361111111, 23754.930555555555, 23754.9375, 23754.944444444445, 23754.95138888889, 23754.958333333332, 23754.965277777777, 23754.972222222223, 23754.979166666668, 23754.98611111111, 23754.993055555555, 23755.0, 23755.006944444445, 23755.01388888889, 23755.020833333332, 23755.027777777777, 23755.034722222223, 23755.041666666668, 23755.04861111111, 23755.055555555555, 23755.0625, 23755.069444444445, 23755.07638888889, 23755.083333333332, 23755.090277777777, 23755.097222222223, 23755.104166666668, 23755.11111111111, 23755.118055555555, 23755.125, 23755.131944444445, 23755.13888888889, 23755.145833333332, 23755.152777777777, 23755.159722222223, 23755.166666666668, 23755.17361111111, 23755.180555555555, 23755.1875, 23755.194444444445, 23755.20138888889, 23755.208333333332, 23755.215277777777, 23755.222222222223, 23755.229166666668, 23755.23611111111, 23755.243055555555, 23755.25, 23755.256944444445, 23755.26388888889, 23755.270833333332, 23755.277777777777, 23755.284722222223, 23755.291666666668, 23755.29861111111, 23755.305555555555, 23755.3125, 23755.319444444445, 23755.32638888889, 23755.333333333332, 23755.340277777777, 23755.347222222223, 23755.354166666668, 23755.36111111111, 23755.368055555555, 23755.375, 23755.381944444445, 23755.38888888889, 23755.395833333332, 23755.402777777777, 23755.409722222223, 23755.416666666668, 23755.42361111111, 23755.430555555555, 23755.4375, 23755.444444444445, 23755.45138888889, 23755.458333333332, 23755.465277777777, 23755.472222222223, 23755.479166666668, 23755.48611111111, 23755.493055555555, 23755.5, 23755.506944444445, 23755.51388888889, 23755.520833333332, 23755.527777777777, 23755.534722222223, 23755.541666666668, 23755.54861111111, 23755.555555555555, 23755.5625, 23755.569444444445, 23755.57638888889, 23755.583333333332, 23755.590277777777, 23755.597222222223, 23755.604166666668, 23755.61111111111, 23755.618055555555, 23755.625, 23755.631944444445, 23755.63888888889, 23755.645833333332, 23755.652777777777, 23755.659722222223, 23755.666666666668, 23755.67361111111, 23755.680555555555, 23755.6875, 23755.694444444445, 23755.70138888889, 23755.708333333332, 23755.715277777777, 23755.722222222223, 23755.729166666668, 23755.73611111111, 23755.743055555555, 23755.75, 23755.756944444445, 23755.76388888889, 23755.770833333332, 23755.777777777777, 23755.784722222223, 23755.791666666668, 23755.79861111111, 23755.805555555555, 23755.8125, 23755.819444444445, 23755.82638888889, 23755.833333333332, 23755.840277777777, 23755.847222222223, 23755.854166666668, 23755.86111111111, 23755.868055555555, 23755.875, 23755.881944444445, 23755.88888888889, 23755.895833333332, 23755.902777777777, 23755.909722222223, 23755.916666666668, 23755.92361111111, 23755.930555555555, 23755.9375, 23755.944444444445, 23755.95138888889, 23755.958333333332, 23755.965277777777, 23755.972222222223, 23755.979166666668, 23755.98611111111, 23755.993055555555, 23756.0, 23756.006944444445, 23756.01388888889, 23756.020833333332, 23756.027777777777, 23756.034722222223, 23756.041666666668, 23756.04861111111, 23756.055555555555, 23756.0625, 23756.069444444445, 23756.07638888889, 23756.083333333332, 23756.090277777777, 23756.097222222223, 23756.104166666668, 23756.11111111111, 23756.118055555555, 23756.125, 23756.131944444445, 23756.13888888889, 23756.145833333332, 23756.152777777777, 23756.159722222223, 23756.166666666668, 23756.17361111111, 23756.180555555555, 23756.1875, 23756.194444444445, 23756.20138888889, 23756.208333333332, 23756.215277777777, 23756.222222222223, 23756.229166666668, 23756.23611111111, 23756.243055555555, 23756.25, 23756.256944444445, 23756.26388888889, 23756.270833333332, 23756.277777777777, 23756.284722222223, 23756.291666666668, 23756.29861111111, 23756.305555555555, 23756.3125, 23756.319444444445, 23756.32638888889, 23756.333333333332, 23756.340277777777, 23756.347222222223, 23756.354166666668, 23756.36111111111, 23756.368055555555, 23756.375, 23756.381944444445, 23756.38888888889, 23756.395833333332, 23756.402777777777, 23756.409722222223, 23756.416666666668, 23756.42361111111, 23756.430555555555, 23756.4375, 23756.444444444445, 23756.45138888889, 23756.458333333332, 23756.465277777777, 23756.472222222223, 23756.479166666668, 23756.48611111111, 23756.493055555555, 23756.5, 23756.506944444445, 23756.51388888889, 23756.520833333332, 23756.527777777777, 23756.534722222223, 23756.541666666668, 23756.54861111111, 23756.555555555555, 23756.5625, 23756.569444444445, 23756.57638888889, 23756.583333333332, 23756.590277777777, 23756.597222222223, 23756.604166666668, 23756.61111111111, 23756.618055555555, 23756.625, 23756.631944444445, 23756.63888888889, 23756.645833333332, 23756.652777777777, 23756.659722222223, 23756.666666666668, 23756.67361111111, 23756.680555555555, 23756.6875, 23756.694444444445, 23756.70138888889, 23756.708333333332, 23756.715277777777, 23756.722222222223, 23756.729166666668, 23756.73611111111, 23756.743055555555, 23756.75, 23756.756944444445, 23756.76388888889, 23756.770833333332, 23756.777777777777, 23756.784722222223, 23756.791666666668, 23756.79861111111, 23756.805555555555, 23756.8125, 23756.819444444445, 23756.82638888889, 23756.833333333332, 23756.840277777777, 23756.847222222223, 23756.854166666668, 23756.86111111111, 23756.868055555555, 23756.875, 23756.881944444445, 23756.88888888889, 23756.895833333332, 23756.902777777777, 23756.909722222223, 23756.916666666668, 23756.92361111111, 23756.930555555555, 23756.9375, 23756.944444444445, 23756.95138888889, 23756.958333333332, 23756.965277777777, 23756.972222222223, 23756.979166666668, 23756.98611111111, 23756.993055555555, 23757.0, 23757.006944444445, 23757.01388888889, 23757.020833333332, 23757.027777777777, 23757.034722222223, 23757.041666666668, 23757.04861111111, 23757.055555555555, 23757.0625, 23757.069444444445, 23757.07638888889, 23757.083333333332, 23757.090277777777, 23757.097222222223, 23757.104166666668, 23757.11111111111, 23757.118055555555, 23757.125, 23757.131944444445, 23757.13888888889, 23757.145833333332, 23757.152777777777, 23757.159722222223, 23757.166666666668, 23757.17361111111, 23757.180555555555, 23757.1875, 23757.194444444445, 23757.20138888889, 23757.208333333332, 23757.215277777777, 23757.222222222223, 23757.229166666668, 23757.23611111111, 23757.243055555555, 23757.25, 23757.256944444445, 23757.26388888889, 23757.270833333332, 23757.277777777777, 23757.284722222223, 23757.291666666668, 23757.29861111111, 23757.305555555555, 23757.3125, 23757.319444444445, 23757.32638888889, 23757.333333333332, 23757.340277777777, 23757.347222222223, 23757.354166666668, 23757.36111111111, 23757.368055555555, 23757.375, 23757.381944444445, 23757.38888888889, 23757.395833333332, 23757.402777777777, 23757.409722222223, 23757.416666666668, 23757.42361111111, 23757.430555555555, 23757.4375, 23757.444444444445, 23757.45138888889, 23757.458333333332, 23757.465277777777, 23757.472222222223, 23757.479166666668, 23757.48611111111, 23757.493055555555, 23757.5, 23757.506944444445, 23757.51388888889, 23757.520833333332, 23757.527777777777, 23757.534722222223, 23757.541666666668, 23757.54861111111, 23757.555555555555, 23757.5625, 23757.569444444445, 23757.57638888889, 23757.583333333332, 23757.590277777777, 23757.597222222223, 23757.604166666668, 23757.61111111111, 23757.618055555555, 23757.625, 23757.631944444445, 23757.63888888889, 23757.645833333332, 23757.652777777777, 23757.659722222223, 23757.666666666668, 23757.67361111111, 23757.680555555555, 23757.6875, 23757.694444444445, 23757.70138888889, 23757.708333333332, 23757.715277777777, 23757.722222222223, 23757.729166666668, 23757.73611111111, 23757.743055555555, 23757.75, 23757.756944444445, 23757.76388888889, 23757.770833333332, 23757.777777777777, 23757.784722222223, 23757.791666666668, 23757.79861111111, 23757.805555555555, 23757.8125, 23757.819444444445, 23757.82638888889, 23757.833333333332, 23757.840277777777, 23757.847222222223, 23757.854166666668, 23757.86111111111, 23757.868055555555, 23757.875, 23757.881944444445, 23757.88888888889, 23757.895833333332, 23757.902777777777, 23757.909722222223, 23757.916666666668, 23757.92361111111, 23757.930555555555, 23757.9375, 23757.944444444445, 23757.95138888889, 23757.958333333332, 23757.965277777777, 23757.972222222223, 23757.979166666668, 23757.98611111111, 23757.993055555555, 23758.0, 23758.006944444445, 23758.01388888889, 23758.020833333332, 23758.027777777777, 23758.034722222223, 23758.041666666668, 23758.04861111111, 23758.055555555555, 23758.0625, 23758.069444444445, 23758.07638888889, 23758.083333333332, 23758.090277777777, 23758.097222222223, 23758.104166666668, 23758.11111111111, 23758.118055555555, 23758.125, 23758.131944444445, 23758.13888888889, 23758.145833333332, 23758.152777777777, 23758.159722222223, 23758.166666666668, 23758.17361111111, 23758.180555555555, 23758.1875, 23758.194444444445, 23758.20138888889, 23758.208333333332, 23758.215277777777, 23758.222222222223, 23758.229166666668, 23758.23611111111, 23758.243055555555, 23758.25, 23758.256944444445, 23758.26388888889, 23758.270833333332, 23758.277777777777, 23758.284722222223, 23758.291666666668, 23758.29861111111, 23758.305555555555, 23758.3125, 23758.319444444445, 23758.32638888889, 23758.333333333332, 23758.340277777777, 23758.347222222223, 23758.354166666668, 23758.36111111111, 23758.368055555555, 23758.375, 23758.381944444445, 23758.38888888889, 23758.395833333332, 23758.402777777777, 23758.409722222223, 23758.416666666668, 23758.42361111111, 23758.430555555555, 23758.4375, 23758.444444444445, 23758.45138888889, 23758.458333333332, 23758.465277777777, 23758.472222222223, 23758.479166666668, 23758.48611111111, 23758.493055555555, 23758.5, 23758.506944444445, 23758.51388888889, 23758.520833333332, 23758.527777777777, 23758.534722222223, 23758.541666666668, 23758.54861111111, 23758.555555555555, 23758.5625, 23758.569444444445, 23758.57638888889, 23758.583333333332, 23758.590277777777, 23758.597222222223, 23758.604166666668, 23758.61111111111, 23758.618055555555, 23758.625, 23758.631944444445, 23758.63888888889, 23758.645833333332, 23758.652777777777, 23758.659722222223, 23758.666666666668, 23758.67361111111, 23758.680555555555, 23758.6875, 23758.694444444445, 23758.70138888889, 23758.708333333332, 23758.715277777777, 23758.722222222223, 23758.729166666668, 23758.73611111111, 23758.743055555555, 23758.75, 23758.756944444445, 23758.76388888889, 23758.770833333332, 23758.777777777777, 23758.784722222223, 23758.791666666668, 23758.79861111111, 23758.805555555555, 23758.8125, 23758.819444444445, 23758.82638888889, 23758.833333333332, 23758.840277777777, 23758.847222222223, 23758.854166666668, 23758.86111111111, 23758.868055555555, 23758.875, 23758.881944444445, 23758.88888888889, 23758.895833333332, 23758.902777777777, 23758.909722222223, 23758.916666666668, 23758.92361111111, 23758.930555555555, 23758.9375, 23758.944444444445, 23758.95138888889, 23758.958333333332, 23758.965277777777, 23758.972222222223, 23758.979166666668, 23758.98611111111, 23758.993055555555, 23759.0, 23759.006944444445, 23759.01388888889, 23759.020833333332, 23759.027777777777, 23759.034722222223, 23759.041666666668, 23759.04861111111, 23759.055555555555, 23759.0625, 23759.069444444445, 23759.07638888889, 23759.083333333332, 23759.090277777777, 23759.097222222223, 23759.104166666668, 23759.11111111111, 23759.118055555555, 23759.125, 23759.131944444445, 23759.13888888889, 23759.145833333332, 23759.152777777777, 23759.159722222223, 23759.166666666668, 23759.17361111111, 23759.180555555555, 23759.1875, 23759.194444444445, 23759.20138888889, 23759.208333333332, 23759.215277777777, 23759.222222222223, 23759.229166666668, 23759.23611111111, 23759.243055555555, 23759.25, 23759.256944444445, 23759.26388888889, 23759.270833333332, 23759.277777777777, 23759.284722222223, 23759.291666666668, 23759.29861111111, 23759.305555555555, 23759.3125, 23759.319444444445, 23759.32638888889, 23759.333333333332, 23759.340277777777, 23759.347222222223, 23759.354166666668, 23759.36111111111, 23759.368055555555, 23759.375, 23759.381944444445, 23759.38888888889, 23759.395833333332, 23759.402777777777, 23759.409722222223, 23759.416666666668, 23759.42361111111, 23759.430555555555, 23759.4375, 23759.444444444445, 23759.45138888889, 23759.458333333332, 23759.465277777777, 23759.472222222223, 23759.479166666668, 23759.48611111111, 23759.493055555555, 23759.5, 23759.506944444445, 23759.51388888889, 23759.520833333332, 23759.527777777777, 23759.534722222223, 23759.541666666668, 23759.54861111111, 23759.555555555555, 23759.5625, 23759.569444444445, 23759.57638888889, 23759.583333333332, 23759.590277777777, 23759.597222222223, 23759.604166666668, 23759.61111111111, 23759.618055555555, 23759.625, 23759.631944444445, 23759.63888888889, 23759.645833333332, 23759.652777777777, 23759.659722222223, 23759.666666666668, 23759.67361111111, 23759.680555555555, 23759.6875, 23759.694444444445, 23759.70138888889, 23759.708333333332, 23759.715277777777, 23759.722222222223, 23759.729166666668, 23759.73611111111, 23759.743055555555, 23759.75, 23759.756944444445, 23759.76388888889, 23759.770833333332, 23759.777777777777, 23759.784722222223, 23759.791666666668, 23759.79861111111, 23759.805555555555, 23759.8125, 23759.819444444445, 23759.82638888889, 23759.833333333332, 23759.840277777777, 23759.847222222223, 23759.854166666668, 23759.86111111111, 23759.868055555555, 23759.875, 23759.881944444445, 23759.88888888889, 23759.895833333332, 23759.902777777777, 23759.909722222223, 23759.916666666668, 23759.92361111111, 23759.930555555555, 23759.9375, 23759.944444444445, 23759.95138888889, 23759.958333333332, 23759.965277777777, 23759.972222222223, 23759.979166666668, 23759.98611111111, 23759.993055555555, 23760.0, 23760.006944444445, 23760.01388888889, 23760.020833333332, 23760.027777777777, 23760.034722222223, 23760.041666666668, 23760.04861111111, 23760.055555555555, 23760.0625, 23760.069444444445, 23760.07638888889, 23760.083333333332, 23760.090277777777, 23760.097222222223, 23760.104166666668, 23760.11111111111, 23760.118055555555, 23760.125, 23760.131944444445, 23760.13888888889, 23760.145833333332, 23760.152777777777, 23760.159722222223, 23760.166666666668, 23760.17361111111, 23760.180555555555, 23760.1875, 23760.194444444445, 23760.20138888889, 23760.208333333332, 23760.215277777777, 23760.222222222223, 23760.229166666668, 23760.23611111111, 23760.243055555555, 23760.25, 23760.256944444445, 23760.26388888889, 23760.270833333332, 23760.277777777777, 23760.284722222223, 23760.291666666668, 23760.29861111111, 23760.305555555555, 23760.3125, 23760.319444444445, 23760.32638888889, 23760.333333333332, 23760.340277777777, 23760.347222222223, 23760.354166666668, 23760.36111111111, 23760.368055555555, 23760.375, 23760.381944444445, 23760.38888888889, 23760.395833333332, 23760.402777777777, 23760.409722222223, 23760.416666666668, 23760.42361111111, 23760.430555555555, 23760.4375, 23760.444444444445, 23760.45138888889, 23760.458333333332, 23760.465277777777, 23760.472222222223, 23760.479166666668, 23760.48611111111, 23760.493055555555, 23760.5, 23760.506944444445, 23760.51388888889, 23760.520833333332, 23760.527777777777, 23760.534722222223, 23760.541666666668, 23760.54861111111, 23760.555555555555, 23760.5625, 23760.569444444445, 23760.57638888889, 23760.583333333332, 23760.590277777777, 23760.597222222223, 23760.604166666668, 23760.61111111111, 23760.618055555555, 23760.625, 23760.631944444445, 23760.63888888889, 23760.645833333332, 23760.652777777777, 23760.659722222223, 23760.666666666668, 23760.67361111111, 23760.680555555555, 23760.6875, 23760.694444444445, 23760.70138888889, 23760.708333333332, 23760.715277777777, 23760.722222222223, 23760.729166666668, 23760.73611111111, 23760.743055555555, 23760.75, 23760.756944444445, 23760.76388888889, 23760.770833333332, 23760.777777777777, 23760.784722222223, 23760.791666666668, 23760.79861111111, 23760.805555555555, 23760.8125, 23760.819444444445, 23760.82638888889, 23760.833333333332, 23760.840277777777, 23760.847222222223, 23760.854166666668, 23760.86111111111, 23760.868055555555, 23760.875, 23760.881944444445, 23760.88888888889, 23760.895833333332, 23760.902777777777, 23760.909722222223, 23760.916666666668, 23760.92361111111, 23760.930555555555, 23760.9375, 23760.944444444445, 23760.95138888889, 23760.958333333332, 23760.965277777777, 23760.972222222223, 23760.979166666668, 23760.98611111111, 23760.993055555555, 23761.0, 23761.006944444445, 23761.01388888889, 23761.020833333332, 23761.027777777777, 23761.034722222223, 23761.041666666668, 23761.04861111111, 23761.055555555555, 23761.0625, 23761.069444444445, 23761.07638888889, 23761.083333333332, 23761.090277777777, 23761.097222222223, 23761.104166666668, 23761.11111111111, 23761.118055555555, 23761.125, 23761.131944444445, 23761.13888888889}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =100.0
TEMP =
  {18.7997, 18.8352, 18.86, 18.9191, 18.9074, 18.8973, 18.9737, 18.9958, 19.0356, 19.0232, 19.0363, 19.0644, 19.0844, 19.1035, 19.1035, 19.0069, 19.1088, 19.2048, 19.0982, 19.1206, 19.0556, 19.06, 19.021, 18.8893, 18.8679, 18.8643, 18.9041, 18.9371, 18.9075, 18.8703, 18.8548, 18.5927, 18.5883, 18.5408, 18.3785, 18.2997, 18.4788, 18.5166, 18.5325, 18.5724, 18.6395, 18.7626, 18.7884, 18.6668, 18.6239, 18.5947, 18.603, 18.5793, 18.4504, 18.4698, 18.5672, 18.5176, 18.5422, 18.4952, 18.4564, 18.498, 18.5687, 18.6035, 18.5868, 18.5272, 18.4944, 18.4846, 18.506, 18.5189, 18.5066, 18.4897, 18.5187, 18.5148, 18.552, 18.5917, 18.6244, 18.6209, 18.7012, 18.727, 18.7381, 18.6733, 18.6545, 18.6979, 18.7062, 18.6689, 18.8062, 18.7334, 18.7795, 18.6342, 18.5736, 18.4592, 18.4484, 18.3478, 18.347, 18.4189, 18.6157, 18.7302, 18.6793, 18.5302, 18.5081, 18.5567, 18.5903, 18.6218, 18.5807, 18.613, 18.65, 18.7184, 18.7066, 18.7257, 18.7086, 18.8507, 18.8004, 18.7918, 18.7368, 18.8449, 18.7565, 18.8365, 18.8305, 18.8303, 18.7918, 18.786, 18.8801, 18.8516, 18.7631, 18.6785, 18.6443, 18.7426, 18.6981, 18.4355, 18.4099, 18.4222, 18.401, 18.3454, 18.3445, 18.2973, 18.3135, 18.4399, 18.3326, 18.312, 18.3039, 18.3188, 18.3762, 18.3981, 18.4174, 18.3939, 18.3703, 18.4235, 18.4568, 18.4437, 18.442, 18.4308, 18.4331, 18.4352, 18.4478, 18.4469, 18.4631, 18.4761, 18.4914, 18.5063, 18.5424, 18.5193, 18.5024, 18.4802, 18.4765, 18.4697, 18.4428, 18.4253, 18.4251, 18.4027, 18.3879, 18.4024, 18.429, 18.422, 18.44, 18.4591, 18.4535, 18.4442, 18.4253, 18.4487, 18.4668, 18.476, 18.4467, 18.4047, 18.3722, 18.3787, 18.4054, 18.3687, 18.3822, 18.4219, 18.397, 18.4015, 18.4117, 18.4168, 18.4584, 18.4709, 18.4783, 18.4834, 18.4839, 18.4719, 18.3767, 18.3812, 18.4811, 18.4947, 18.493, 18.4954, 18.4873, 18.4897, 18.4893, 18.4883, 18.451, 18.4355, 18.4581, 18.4579, 18.4466, 18.4565, 18.4647, 18.4771, 18.4829, 18.498, 18.6252, 18.6902, 18.4677, 18.4452, 18.4346, 18.4914, 18.4709, 18.4286, 18.5278, 18.5682, 18.5591, 18.5758, 18.4812, 18.5708, 18.6033, 18.6315, 18.7028, 18.7811, 18.8582, 18.773, 18.8422, 18.7806, 18.878, 18.9483, 18.8769, 18.7505, 18.7784, 18.6771, 18.6356, 18.5008, 18.4021, 18.3867, 18.3896, 18.4002, 18.394, 18.3829, 18.3782, 18.4077, 18.3795, 18.3254, 18.325, 18.3075, 18.2949, 18.2812, 18.3, 18.2901, 18.29, 18.3011, 18.3072, 18.2869, 18.2929, 18.3011, 18.3104, 18.2977, 18.2709, 18.2626, 18.2639, 18.2631, 18.2643, 18.2675, 18.2654, 18.2671, 18.2687, 18.2711, 18.2739, 18.266, 18.2803, 18.3312, 18.2821, 18.2752, 18.2708, 18.2709, 18.2766, 18.278, 18.2764, 18.2824, 18.2813, 18.284, 18.2785, 18.2801, 18.2768, 18.2042, 18.2375, 18.2573, 18.2649, 18.2209, 18.2084, 18.1963, 18.1764, 18.1978, 18.2415, 18.2576, 18.2545, 18.2447, 18.2475, 18.2693, 18.2848, 18.3714, 18.3011, 18.2901, 18.2986, 18.4719, 18.4686, 18.7842, 18.7746, 18.495, 18.4311, 18.4595, 18.4985, 18.3189, 18.3279, 18.3253, 18.2699, 18.334, 18.4944, 18.4587, 18.7986, 18.594, 18.7123, 18.7901, 18.5252, 18.4322, 18.3521, 18.3499, 18.3831, 18.4279, 18.5521, 18.4946, 18.5877, 18.4397, 18.4148, 18.3758, 18.3504, 18.3787, 18.3704, 18.3934, 18.4199, 18.4933, 18.5172, 18.4951, 18.411, 18.3577, 18.2648, 18.3379, 18.2769, 18.3269, 18.2548, 18.2861, 18.3005, 18.2248, 18.207, 18.2064, 18.3439, 18.3917, 18.3425, 18.321, 18.3741, 18.377, 18.3757, 18.387, 18.3965, 18.3816, 18.3948, 18.4005, 18.4133, 18.4263, 18.4196, 18.4438, 18.4103, 18.4384, 18.422, 18.4255, 18.4431, 18.4034, 18.4164, 18.4205, 18.3734, 18.3333, 18.204, 18.2058, 18.2085, 18.0856, 18.0552, 18.0039, 17.9933, 18.0459, 18.0081, 18.2402, 18.2521, 18.3004, 18.2578, 18.2661, 18.0034, 18.2054, 18.2696, 18.3564, 18.303, 18.2753, 18.1574, 18.2048, 18.1603, 18.1733, 18.3443, 18.2766, 18.3586, 18.2079, 18.1201, 18.1422, 18.1607, 18.107, 18.1101, 18.107, 18.0542, 18.0448, 18.0521, 18.1122, 18.1666, 18.0739, 18.1068, 18.3522, 18.156, 18.2126, 18.2129, 18.2985, 18.1021, 18.0759, 18.0547, 18.0314, 18.021, 17.9529, 18.0103, 18.0058, 18.1373, 18.059, 18.0273, 18.0268, 17.9973, 18.0823, 18.167, 18.2173, 18.2274, 18.1948, 18.1854, 18.1388, 18.1518, 18.1725, 18.195, 18.1551, 18.1346, 18.1271, 18.1772, 18.183, 18.2102, 18.208, 18.1706, 18.2112, 18.2126, 18.2213, 18.2134, 18.1624, 18.1554, 18.1428, 18.1593, 18.2876, 18.2877, 18.2861, 18.2391, 18.2574, 18.3298, 18.3514, 18.3184, 18.2724, 18.2599, 18.2873, 18.2643, 18.2768, 18.3042, 18.3093, 18.2849, 18.2712, 18.2835, 18.3004, 18.2516, 18.2535, 18.2472, 18.239, 18.2458, 18.2278, 18.2197, 18.2108, 18.4485, 18.2105, 18.2985, 18.2133, 18.4451, 18.4166, 18.5448, 18.4901, 18.4267, 18.3576, 18.2263, 18.436, 18.3944, 18.5096, 18.5176, 18.4658, 18.446, 18.5071, 18.471, 18.5044, 18.4916, 18.4766, 18.5002, 18.5005, 18.5262, 18.6089, 18.5087, 18.4262, 18.4187, 18.4344, 18.4701, 18.468, 18.4425, 18.2418, 18.3571, 18.2608, 18.2055, 18.1732, 18.139, 18.2694, 18.0531, 18.0541, 18.0299, 18.0612, 18.2825, 18.4704, 18.4547, 18.3643, 18.1238, 17.9149, 17.8365, 17.8569, 18.1005, 18.1722, 18.1271, 18.0862, 18.1039, 18.1992, 18.2055, 18.1573, 18.1303, 18.0671, 18.0723, 18.067, 18.0753, 18.0899, 18.0407, 18.1065, 18.108, 18.0471, 18.0493, 18.0494, 18.0202, 18.0228, 18.0421, 18.0539, 17.9888, 17.9867, 17.9572, 17.953, 17.9386, 17.9349, 17.8528, 17.9387, 17.9965, 18.0632, 18.0269, 18.0735, 18.0334, 18.0182, 18.0291, 18.0316, 18.0694, 18.0692, 18.0757, 18.071, 18.154, 18.1772, 18.1836, 18.1293, 18.1245, 18.1949, 18.1916, 18.1879, 18.1873, 18.1737, 18.1767, 18.187, 18.1827, 18.1988, 18.2034, 18.2, 18.2046, 18.218, 18.2311, 18.2338, 18.2392, 18.2433, 18.2445, 18.2482, 18.1527, 18.1767, 18.1595, 18.1711, 18.2544, 18.2581, 18.2612, 18.2397, 18.1674, 18.2542, 18.1446, 18.1414, 18.1428, 18.1464, 18.166, 18.184, 18.1613, 18.1874, 18.245, 18.2451, 18.2231, 18.2007, 18.245, 18.2472, 18.2777, 18.2924, 18.2959, 18.3039, 18.3139, 18.3089, 18.3077, 18.3065, 18.3128, 18.321, 18.3037, 18.2721, 18.2929, 18.33, 18.2554, 18.3537, 18.5761, 18.3623, 18.4941, 18.3721, 18.4333, 18.276, 18.3775, 18.3624, 18.3585, 18.5083, 18.352, 18.2776, 18.2765, 18.2873, 18.281, 18.2553, 18.1959, 18.2711, 18.2128, 18.1922, 18.1754, 18.197, 18.2266, 18.2286, 18.1792, 18.1684, 18.1595, 18.1477, 18.1467, 18.2945, 18.132, 18.1118, 18.1082, 18.0915, 18.0227, 17.9825, 17.9681, 17.9555, 17.9488, 17.9444, 17.9338, 17.9186, 17.954, 18.0919, 18.1307, 18.0883, 18.0762, 18.0759, 18.0804, 18.0707, 18.0943, 18.0987, 18.1015, 18.0422, 18.0628, 18.0597, 18.0537, 18.0499, 17.9225, 17.8998, 17.9316, 17.9658, 17.9856, 18.017, 18.0293, 17.9621, 17.8911, 17.9434, 17.9996, 17.9562, 17.9314, 17.9135, 17.8799, 17.8299, 17.7922, 17.815, 17.8774, 17.9197, 17.8542, 17.9318, 17.9605, 18.0633, 18.0, 18.0622, 18.0548, 18.1216, 18.2067, 18.2225, 18.2228, 18.2343, 18.1953, 18.1953, 18.2499, 18.1577, 18.0167, 18.0067, 17.9743, 17.9957, 18.0126, 18.0357, 18.0275, 17.9508, 18.0119, 18.0237, 18.0484, 18.0733, 18.0306, 18.1607, 18.1054, 18.1221, 17.9906, 18.0669, 17.9941, 17.9933, 18.1364, 18.0252, 18.2657, 18.3051, 18.2949, 18.3477, 18.3379, 18.3176, 18.2841, 18.2401, 18.1719, 18.2909, 18.2681, 18.3109, 18.3027, 18.4061, 18.2347, 18.3371, 18.2258, 18.2206, 18.2158, 18.3446, 18.1798, 18.1599, 18.3396, 18.1586, 18.0626, 18.0231, 18.0209, 18.0286, 17.9998, 17.9859, 17.9927, 18.1902, 18.1315, 18.0174, 18.067, 18.0539, 18.1829, 18.1308, 18.2074, 18.1714, 18.2528, 18.1939, 18.2634, 18.321, 18.1993, 18.2059, 18.2019, 18.2848, 18.4533, 18.3938, 18.2886, 18.4395, 18.286, 18.3433, 18.221, 18.2083, 18.1649, 18.1688, 18.2097, 18.1554, 18.2584, 18.2305, 18.2297, 18.3115, 18.2463, 18.2926, 18.1449, 18.1349, 18.3572, 18.1715, 17.9886, 18.1542, 18.2119, 18.1549, 18.1596, 18.3227, 18.1099, 18.1489, 18.183, 18.1687, 18.1633, 18.1439, 18.1272, 18.1071, 18.1145, 18.2334, 18.2205, 18.2349, 18.1573, 18.0643, 18.147, 18.0242, 18.071, 18.0758, 18.0319, 18.0488, 17.993, 17.9771, 17.9682, 17.9749, 17.9418, 17.9234, 17.9252, 17.9102, 17.8756, 17.8671, 17.8592, 21.4047, 23.8757, 23.0044, 23.8901, 23.8627, 23.7329, 22.9613, 22.3277, 22.0586, 22.0005, 22.1319, 22.1067, 22.1921, 22.2597, 22.3604, 22.649, 24.5655, 25.5712, 26.4362, 27.6535, 28.1111, 27.9759, 27.8995, 27.818, 27.7648, 27.7292, 27.6791, 27.629, 27.5671, 27.5012, 27.4343, 27.3642, 27.2903, 27.2073, 27.1326, 27.0528, 26.9732, 26.8991, 26.8263, 26.757, 26.6788, 26.5947, 26.5181, 26.4438, 26.3798, 26.31, 26.2424, 26.1738, 26.0977, 26.0268, 25.9539, 25.8798, 25.8074, 25.728, 25.6452, 25.5537, 25.4751, 25.3903, 25.3108, 25.2354, 25.1672, 25.0921, 25.0196, 24.9484, 24.8803, 24.8152, 24.7523, 24.6936, 24.6341, 24.5764, 24.5211, 24.4642, 24.4115, 24.3553, 24.2997, 24.2429, 24.1824, 24.1123, 24.0443, 23.9761, 23.9066, 23.8207, 23.7447, 23.6681, 23.5995, 23.5413, 23.4894, 23.4449, 23.4032, 23.3661, 23.3301, 23.2912, 23.2438, 23.192, 23.1336, 23.075, 23.0222, 22.9608, 22.9035, 22.843, 22.7858, 22.7271, 22.6661, 22.5997, 22.5464, 22.4833, 22.4302, 22.3751, 22.3196, 22.2609, 22.2073, 22.1545, 22.0916, 22.0364, 21.9822, 21.9245, 21.8695, 21.8184, 21.7693, 21.7254, 21.681, 21.64, 21.6024, 21.57, 21.5357, 21.5062, 21.479, 21.4527, 21.4312, 21.4117, 21.3914, 21.3739, 21.3582, 21.3442, 21.3391, 21.3359, 21.3315, 21.3292, 21.3272, 21.3272, 21.3377, 21.3549, 21.3629, 21.3679, 21.3771, 21.3872, 21.3977, 21.409}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_REL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
DEPTH =
  {110.919205, 110.70322, 110.73091, 110.75643, 110.83077, 110.77794, 110.76826, 110.77428, 110.710014, 110.74564, 110.89494, 110.74704, 110.72395, 110.87171, 110.6912, 110.86417, 110.80846, 110.697845, 110.87156, 110.84222, 110.71328, 110.92288, 110.87763, 110.91729, 110.93818, 110.95805, 110.89044, 110.77334, 110.87393, 110.82139, 110.84936, 110.79348, 110.87395, 110.917816, 110.96475, 110.9455, 111.000046, 111.00777, 110.958145, 110.95824, 110.94747, 111.05741, 111.00829, 110.88133, 111.0421, 110.94364, 110.973526, 110.94238, 111.00255, 110.89867, 111.039505, 111.03107, 111.06173, 111.103806, 110.98432, 111.04834, 110.94933, 110.890625, 111.030685, 111.01447, 110.94564, 110.96019, 111.09022, 111.027245, 110.983826, 111.09581, 110.97125, 110.98978, 111.00685, 110.98647, 111.04299, 111.01483, 111.04678, 111.096375, 111.0419, 111.09207, 111.080475, 110.896324, 111.05904, 110.99858, 110.94094, 110.916824, 111.04452, 111.017204, 110.88524, 111.029625, 110.87996, 110.96007, 110.91336, 110.94729, 110.89442, 110.95075, 110.97684, 110.95438, 110.98642, 110.89323, 110.8146, 110.84798, 110.800354, 110.76305, 110.77316, 110.77684, 110.858475, 110.72298, 110.67218, 110.895195, 110.74832, 110.82797, 110.74556, 110.76732, 110.8071, 110.864746, 110.89273, 110.78397, 110.770035, 110.7449, 110.7563, 110.67179, 110.67204, 110.714294, 110.694, 110.71423, 110.674324, 110.71389, 110.60852, 110.68187, 110.6113, 110.71196, 110.73931, 110.57075, 110.74007, 110.60294, 110.74628, 110.68347, 110.55857, 110.55532, 110.58382, 110.51332, 110.66199, 110.63165, 110.535095, 110.66017, 110.58562, 110.63235, 110.65329, 110.668144, 110.575035, 110.66138, 110.60921, 110.71732, 110.7776, 110.699814, 110.69084, 110.66698, 110.71343, 110.62137, 110.693565, 110.70233, 110.72435, 110.708595, 110.76622, 110.76275, 110.835686, 110.732925, 110.788086, 110.67574, 110.77027, 110.79641, 110.8836, 110.731926, 110.76837, 110.80269, 110.81591, 110.84496, 110.74214, 110.86383, 110.806244, 110.73429, 110.729225, 110.81071, 110.971466, 110.87191, 110.85298, 110.96594, 110.86482, 110.822174, 110.90715, 110.9594, 110.86144, 110.87549, 110.80274, 110.949585, 110.998344, 110.893036, 110.90713, 110.980064, 110.94448, 110.933266, 111.022934, 110.980896, 111.04591, 110.95082, 110.9257, 111.068214, 111.039795, 111.01852, 110.96894, 110.94942, 111.03453, 111.060616, 111.03269, 110.94958, 111.04303, 111.07688, 110.96637, 111.02168, 110.94534, 111.08732, 110.944214, 111.00154, 111.005646, 110.9763, 110.877914, 110.90476, 110.91822, 110.93339, 110.87846, 110.96826, 110.9662, 110.87955, 110.89861, 110.822624, 111.03428, 110.77311, 110.93414, 110.89149, 110.820404, 110.845566, 110.82771, 110.81008, 110.75455, 110.7379, 110.6759, 110.782135, 110.75124, 110.64895, 110.6512, 110.66694, 110.70762, 110.64341, 110.84754, 110.685936, 110.58012, 110.606384, 110.78061, 110.674904, 110.4872, 110.58166, 110.72171, 110.60077, 110.6932, 110.60773, 110.67124, 110.51753, 110.578865, 110.52493, 110.551895, 110.60884, 110.56507, 110.59056, 110.547745, 110.67247, 110.62508, 110.62915, 110.58438, 110.66966, 110.56197, 110.72775, 110.53805, 110.44248, 110.6207, 110.607864, 110.63989, 110.5372, 110.60511, 110.594536, 110.574585, 110.62451, 110.62982, 110.74959, 110.58747, 110.61432, 110.63939, 110.698074, 110.63516, 110.64514, 110.71243, 110.64084, 110.67544, 110.78725, 110.69127, 110.62552, 110.71295, 110.81146, 110.82089, 110.74095, 110.74234, 110.85799, 110.78823, 110.75921, 110.75867, 110.866646, 110.7191, 110.56322, 110.75978, 110.83078, 110.844185, 110.76583, 110.85018, 110.789185, 110.77619, 110.96659, 110.93431, 110.73668, 110.88313, 110.89459, 110.79146, 110.93035, 110.90674, 110.80687, 110.952065, 110.94469, 110.903564, 111.009514, 110.97551, 110.90827, 110.978424, 110.940414, 111.029655, 111.01714, 111.11284, 111.03596, 111.12967, 111.0647, 111.06472, 111.00002, 111.12675, 111.13363, 111.14224, 111.15867, 111.06328, 111.161446, 111.11027, 111.18532, 110.99756, 111.10972, 111.12879, 111.11002, 111.03305, 111.03398, 111.0571, 111.17115, 111.11995, 111.193016, 111.21155, 110.95362, 110.991745, 111.01276, 111.191444, 111.01141, 110.9738, 111.03536, 111.04813, 110.978874, 111.029045, 110.99543, 111.16219, 111.06033, 110.88753, 110.95934, 110.939674, 110.89165, 110.85179, 110.90662, 110.78639, 110.897125, 110.8402, 110.89756, 110.76601, 110.8126, 110.78051, 110.806854, 110.62271, 110.81824, 110.73507, 110.668625, 110.685776, 110.703514, 110.77, 110.676315, 110.62419, 110.70861, 110.50443, 110.62614, 110.62456, 110.49608, 110.41284, 110.66606, 110.61964, 110.54012, 110.44443, 110.67142, 110.45671, 110.47195, 110.63666, 110.71319, 110.64977, 110.5783, 110.469696, 110.641, 110.61887, 110.52449, 110.49432, 110.6125, 110.51492, 110.55223, 110.65376, 110.54491, 110.63463, 110.577286, 110.577774, 110.45236, 110.534134, 110.65041, 110.58365, 110.60609, 110.654465, 110.612625, 110.58465, 110.57598, 110.59816, 110.76321, 110.73246, 110.647385, 110.75016, 110.752014, 110.67111, 110.73938, 110.74667, 110.7408, 110.82139, 110.73336, 110.83083, 110.78818, 110.73527, 110.85135, 110.80573, 110.785286, 110.83757, 110.94455, 110.79296, 110.890884, 110.82384, 110.95001, 110.71724, 110.94719, 110.779495, 110.91491, 110.847946, 110.880585, 110.82386, 110.805016, 110.9155, 110.92258, 111.062775, 111.0105, 110.91808, 110.933235, 110.97616, 110.89023, 110.980865, 110.91635, 111.08946, 111.13167, 111.02633, 111.053535, 111.13195, 111.24069, 111.166565, 111.01874, 111.028885, 111.13356, 111.2387, 111.21046, 111.19272, 111.05837, 111.09898, 111.23094, 111.19715, 111.36661, 111.18512, 111.196686, 111.37032, 111.1937, 111.14961, 111.29118, 111.31693, 111.15994, 111.21836, 111.10849, 111.229355, 111.22036, 111.17517, 111.14761, 111.234665, 111.152916, 111.067635, 111.08224, 111.225334, 111.05634, 111.19243, 111.22192, 111.04966, 111.12969, 111.05466, 110.9256, 110.993484, 111.093216, 110.84768, 110.91499, 110.91066, 110.81369, 110.89799, 110.837296, 110.86825, 110.80132, 110.838394, 110.79862, 110.72356, 110.83923, 110.748566, 110.7626, 110.62118, 110.647255, 110.52444, 110.74782, 110.51323, 110.58565, 110.52958, 110.61451, 110.52348, 110.38318, 110.55288, 110.75597, 110.58131, 110.445915, 110.62285, 110.51797, 110.5988, 110.53157, 110.51091, 110.60059, 110.41678, 110.52859, 110.67433, 110.43995, 110.57097, 110.61805, 110.466995, 110.61304, 110.64246, 110.60636, 110.64418, 110.44, 110.4494, 110.51977, 110.60749, 110.653, 110.574135, 110.6358, 110.6996, 110.73047, 110.68729, 110.673416, 110.68288, 110.63407, 110.70593, 110.80232, 110.821396, 110.89369, 110.914345, 110.85756, 110.89207, 110.7839, 110.73651, 110.85397, 110.90332, 110.744026, 110.86809, 110.985, 110.816696, 110.89135, 110.76724, 110.904465, 110.79119, 110.84071, 110.70996, 110.85088, 110.89817, 110.91757, 110.808655, 110.85028, 110.864716, 110.83011, 110.96101, 111.05397, 111.129005, 110.95443, 111.054504, 110.97883, 111.01818, 110.99484, 111.05856, 110.904205, 111.00499, 110.866646, 111.04786, 110.96887, 111.208664, 111.02072, 111.04027, 111.07457, 111.03702, 111.10586, 111.00989, 111.01766, 111.03548, 111.1262, 111.13922, 111.05119, 111.19226, 111.11368, 111.22965, 111.059296, 111.19127, 111.16801, 111.22096, 111.18784, 111.31008, 111.23191, 111.24223, 111.17599, 111.1638, 111.20581, 111.261406, 111.26146, 111.093185, 111.173775, 111.190125, 111.127785, 111.15979, 111.21987, 111.14778, 111.27944, 111.19614, 111.11641, 111.17821, 111.172195, 111.158615, 111.12485, 110.99428, 110.98172, 111.08494, 110.87717, 110.94091, 110.94081, 111.0029, 110.98776, 110.806274, 110.778305, 110.88016, 110.857285, 110.763954, 111.03407, 110.76188, 110.76493, 110.66651, 110.64424, 110.72764, 110.60618, 110.54161, 110.66778, 110.660675, 110.63711, 110.634964, 110.59364, 110.545975, 110.52803, 110.5359, 110.6484, 110.53186, 110.4802, 110.46338, 110.48581, 110.49007, 110.5349, 110.55323, 110.53438, 110.42746, 110.496445, 110.41228, 110.46204, 110.65977, 110.45549, 110.47197, 110.39409, 110.400375, 110.40957, 110.64856, 110.66601, 110.59884, 110.51783, 110.49715, 110.68208, 110.57036, 110.75825, 110.599655, 110.58328, 110.70124, 110.69386, 110.5381, 110.70041, 110.575424, 110.738815, 110.702675, 110.7337, 110.74351, 110.81697, 110.798676, 110.77635, 110.65482, 110.82124, 110.73135, 110.77323, 110.80237, 110.73475, 110.78894, 110.804825, 110.72837, 110.851, 110.78611, 110.7931, 110.75694, 110.68495, 110.75014, 110.79766, 110.85285, 110.821304, 110.75808, 110.77026, 110.84062, 110.837326, 110.82358, 110.906586, 110.885826, 110.80443, 110.874115, 110.92472, 110.94583, 110.90164, 110.86795, 110.8985, 110.982666, 110.91954, 110.95311, 110.97215, 110.948074, 111.01594, 111.047165, 110.97954, 111.01678, 111.035324, 111.04378, 111.10606, 111.0634, 111.0708, 111.118286, 111.1816, 111.15177, 111.30859, 111.08542, 111.31881, 111.18783, 111.30028, 111.1608, 111.21406, 111.20098, 111.26576, 111.17163, 111.23616, 111.24667, 111.289444, 111.33174, 111.27092, 111.285225, 111.29736, 111.22183, 111.3593, 111.15935, 111.284225, 111.26138, 111.303604, 111.2397, 111.201836, 111.292206, 111.32179, 111.25978, 110.99218, 111.220825, 111.03572, 111.15297, 111.005035, 111.07998, 111.00412, 110.91668, 111.01657, 110.94903, 110.90858, 110.972, 110.83442, 110.86172, 110.94517, 110.804115, 110.83741, 110.879944, 110.756226, 110.80754, 110.70359, 110.72316, 110.64316, 110.71518, 110.52066, 110.580376, 110.70415, 110.69001, 110.66224, 110.641106, 110.53654, 110.59598, 110.53956, 110.5878, 110.5786, 110.529625, 110.55091, 110.61362, 110.605484, 110.50927, 110.60441, 110.59848, 110.73656, 110.60057, 110.69411, 110.669914, 110.57438, 110.63942, 110.72763, 110.75, 110.83876, 110.69939, 110.65086, 110.88979, 110.707886, 110.7082, 110.917114, 110.79167, 110.84784, 110.8343, 110.92095, 110.951744, 111.04355, 110.98429, 111.09146, 110.94043, 111.193405, 110.95178, 111.03894, 109.27545, 33.8999, 1.6033775, 0.14835767, 0.12171414, 0.11795545, 0.118888594, 0.18825305, 0.12337086, 0.12010125, 0.11926668, 0.12079117, 0.11389377, 0.11745907, 0.113193884, 0.107979, 0.107151404, 0.10549096, 0.09585886, 0.08759834, 0.0703091, 0.19602352, 0.1813009, 0.17385778, 0.20599665, 0.20931861, 0.20710945, 0.20489341, 0.20062375, 0.20213045, 0.19897863, 0.19580099, 0.19786191, 0.19731289, 0.19648068, 0.19015191, 0.19070384, 0.19097888, 0.18837433, 0.19043222, 0.18781427, 0.19098619, 0.1878112, 0.18836129, 0.19263971, 0.19208342, 0.1920819, 0.19524202, 0.1984138, 0.19664365, 0.19774306, 0.19717678, 0.19746435, 0.20118734, 0.19912338, 0.20462021, 0.20461388, 0.20310287, 0.20655683, 0.20709956, 0.20560059, 0.208216, 0.20710626, 0.20504096, 0.20820305, 0.2087587, 0.2098676, 0.21014383, 0.20960152, 0.21069634, 0.21153322, 0.21469218, 0.21153545, 0.21154101, 0.20947874, 0.21208224, 0.21208356, 0.21208054, 0.21580139, 0.21402851, 0.2171885, 0.2177484, 0.21774112, 0.21716963, 0.21979046, 0.2203508, 0.22406942, 0.22091067, 0.22090587, 0.2188504, 0.21996224, 0.22256897, 0.22146136, 0.2168043, 0.22023183, 0.2213515, 0.2213515, 0.21846123, 0.2178983, 0.21995074, 0.2173426, 0.22050473, 0.2173426, 0.22022697, 0.22133812, 0.22245428, 0.22822219, 0.22822785, 0.22878426, 0.22671792, 0.2324837, 0.23193383, 0.22958925, 0.23070583, 0.23125449, 0.23153222, 0.2315391, 0.23097369, 0.23415048, 0.23842907, 0.2346985, 0.23441333, 0.23496577, 0.23496155, 0.23551753, 0.23661959, 0.24183637, 0.23978812, 0.24348944, 0.24611461, 0.24322876, 0.24527678, 0.24267021, 0.24294558, 0.24350931, 0.24611199, 0.24583815, 0.24267904, 0.24267164, 0.24294984, 0.24872273, 0.24555111, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
