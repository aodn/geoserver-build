netcdf file-120.nc {
  dimensions:
    DEPTH = 20;
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593, 22988.062905092593}
TEMP =
  {32.0631, 32.0617, 32.0501, 32.0083, 31.9795, 31.9654, 31.9528, 31.94, 31.9295, 31.9192, 31.9059, 31.8936, 31.8871, 31.8838, 31.879, 31.8777, 31.8747, 31.8657, 31.8641, 31.8636}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879, 21.873}
}
