netcdf file-115.nc {
  dimensions:
    DEPTH = 20;
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889, 22987.85763888889}
TEMP =
  {31.8454, 31.9199, 31.9188, 31.9228, 31.9237, 31.9227, 31.9208, 31.9232, 31.9236, 31.9246, 31.9235, 31.9231, 31.9244, 31.925, 31.9263, 31.9275, 31.9278, 31.9283, 31.9286, 31.9283}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89, 19.884, 20.878}
}
