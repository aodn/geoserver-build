netcdf file-108.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (20 currently)
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926, 22659.27207175926}
TEMP =
  {31.5306, 31.5328, 31.5345, 31.5317, 31.5314, 31.5308, 31.5298, 31.5308, 31.5307, 31.5301, 31.5277, 31.519, 31.5154, 31.5138, 31.5131, 31.5124, 31.5133, 31.5142, 31.5137, 31.5138}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.891, 19.885}
}
