netcdf file-96.nc {
  dimensions:
    DEPTH = 21;
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445, 22658.772256944445}
TEMP =
  {31.5209, 31.5237, 31.5287, 31.5278, 31.5302, 31.5346, 31.5366, 31.5389, 31.5405, 31.5416, 31.5425, 31.544, 31.5454, 31.5458, 31.5452, 31.5443, 31.5436, 31.5434, 31.5436, 31.5424, 31.5413}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89, 19.885, 20.879}
}
