netcdf file-58.nc {
  dimensions:
    DEPTH = 48;
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407, 23123.128032407407}
TEMP =
  {22.9263, 22.9269, 22.9252, 22.9244, 22.9229, 22.9165, 22.9131, 22.9121, 22.9106, 22.9095, 22.9078, 22.9062, 22.9047, 22.9039, 22.9027, 22.8997, 22.8979, 22.8967, 22.8949, 22.8923, 22.8911, 22.8903, 22.8908, 22.8916, 22.893, 22.8941, 22.8991, 22.9029, 22.9045, 22.9047, 22.9023, 22.8833, 22.8474, 22.8129, 22.7852, 22.7657, 22.7365, 22.6948, 22.6743, 22.6729, 22.6674, 22.6622, 22.6571, 22.657, 22.6555, 22.6558, 22.6565, 22.6565}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
