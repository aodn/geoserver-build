netcdf file-173.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (26 currently)
  variables:
    float LATITUDE(DEPTH=26);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=26);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=26);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=26);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=26);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=26);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148, 22811.03616898148}
TEMP =
  {22.916, 22.9155, 22.9161, 22.9137, 22.9087, 22.9065, 22.9067, 22.9048, 22.9011, 22.9, 22.9, 22.8978, 22.8977, 22.8957, 22.8948, 22.8953, 22.8957, 22.8946, 22.8943, 22.8943, 22.8945, 22.8946, 22.8946, 22.8943, 22.8942, 22.8947}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835}
}
