netcdf IMOS_ANMN-TS_20150113T230001Z_WATR20_FV01_WATR20-1407-Seabird-SBE37-SM-2000m-P-70_END-20150121T050001Z_id-7739.nc {
  dimensions:
    TIME = 1045;
  variables:
    double TIME(TIME=1045);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=1045);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=1045);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=1045);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=1045);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=1045);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=1045);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=1045);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=1045);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=1045);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=1045);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=1045);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=1045);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been filled using the DEPTH median (mooring).";
  :instrument = "Seabird SBE37-SM (2000m + P)";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "10030";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 70.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = -0.068f; // float
  :geospatial_vertical_max = 81.141f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:01Z";
  :time_coverage_end = "2015-01-21T05:00:01Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.95834490741, 23753.96528935185, 23753.972233796296, 23753.97917824074, 23753.986122685186, 23753.993067129628, 23754.000011574073, 23754.00695601852, 23754.013900462964, 23754.02084490741, 23754.02778935185, 23754.034733796296, 23754.04167824074, 23754.048622685186, 23754.055567129628, 23754.062511574073, 23754.06945601852, 23754.076400462964, 23754.08334490741, 23754.09028935185, 23754.097233796296, 23754.10417824074, 23754.111122685186, 23754.118067129628, 23754.125011574073, 23754.13195601852, 23754.138900462964, 23754.14584490741, 23754.15278935185, 23754.159733796296, 23754.16667824074, 23754.173622685186, 23754.180567129628, 23754.187511574073, 23754.19445601852, 23754.201400462964, 23754.20834490741, 23754.21528935185, 23754.222233796296, 23754.22917824074, 23754.236122685186, 23754.243067129628, 23754.250011574073, 23754.25695601852, 23754.263900462964, 23754.27084490741, 23754.27778935185, 23754.284733796296, 23754.29167824074, 23754.298622685186, 23754.305567129628, 23754.312511574073, 23754.31945601852, 23754.326400462964, 23754.33334490741, 23754.34028935185, 23754.347233796296, 23754.35417824074, 23754.361122685186, 23754.368067129628, 23754.375011574073, 23754.38195601852, 23754.388900462964, 23754.39584490741, 23754.40278935185, 23754.409733796296, 23754.41667824074, 23754.423622685186, 23754.430567129628, 23754.437511574073, 23754.44445601852, 23754.451400462964, 23754.45834490741, 23754.46528935185, 23754.472233796296, 23754.47917824074, 23754.486122685186, 23754.493067129628, 23754.500011574073, 23754.50695601852, 23754.513900462964, 23754.52084490741, 23754.52778935185, 23754.534733796296, 23754.54167824074, 23754.548622685186, 23754.555567129628, 23754.562511574073, 23754.56945601852, 23754.576400462964, 23754.58334490741, 23754.59028935185, 23754.597233796296, 23754.60417824074, 23754.611122685186, 23754.618067129628, 23754.625011574073, 23754.63195601852, 23754.638900462964, 23754.64584490741, 23754.65278935185, 23754.659733796296, 23754.66667824074, 23754.673622685186, 23754.680567129628, 23754.687511574073, 23754.69445601852, 23754.701400462964, 23754.70834490741, 23754.71528935185, 23754.722233796296, 23754.72917824074, 23754.736122685186, 23754.743067129628, 23754.750011574073, 23754.75695601852, 23754.763900462964, 23754.77084490741, 23754.77778935185, 23754.784733796296, 23754.79167824074, 23754.798622685186, 23754.805567129628, 23754.812511574073, 23754.81945601852, 23754.826400462964, 23754.83334490741, 23754.84028935185, 23754.847233796296, 23754.85417824074, 23754.861122685186, 23754.868067129628, 23754.875011574073, 23754.88195601852, 23754.888900462964, 23754.89584490741, 23754.90278935185, 23754.909733796296, 23754.91667824074, 23754.923622685186, 23754.930567129628, 23754.937511574073, 23754.94445601852, 23754.951400462964, 23754.95834490741, 23754.96528935185, 23754.972233796296, 23754.97917824074, 23754.986122685186, 23754.993067129628, 23755.000011574073, 23755.00695601852, 23755.013900462964, 23755.02084490741, 23755.02778935185, 23755.034733796296, 23755.04167824074, 23755.048622685186, 23755.055567129628, 23755.062511574073, 23755.06945601852, 23755.076400462964, 23755.08334490741, 23755.09028935185, 23755.097233796296, 23755.10417824074, 23755.111122685186, 23755.118067129628, 23755.125011574073, 23755.13195601852, 23755.138900462964, 23755.14584490741, 23755.15278935185, 23755.159733796296, 23755.16667824074, 23755.173622685186, 23755.180567129628, 23755.187511574073, 23755.19445601852, 23755.201400462964, 23755.20834490741, 23755.21528935185, 23755.222233796296, 23755.22917824074, 23755.236122685186, 23755.243067129628, 23755.250011574073, 23755.25695601852, 23755.263900462964, 23755.27084490741, 23755.27778935185, 23755.284733796296, 23755.29167824074, 23755.298622685186, 23755.305567129628, 23755.312511574073, 23755.31945601852, 23755.326400462964, 23755.33334490741, 23755.34028935185, 23755.347233796296, 23755.35417824074, 23755.361122685186, 23755.368067129628, 23755.375011574073, 23755.38195601852, 23755.388900462964, 23755.39584490741, 23755.40278935185, 23755.409733796296, 23755.41667824074, 23755.423622685186, 23755.430567129628, 23755.437511574073, 23755.44445601852, 23755.451400462964, 23755.45834490741, 23755.46528935185, 23755.472233796296, 23755.47917824074, 23755.486122685186, 23755.493067129628, 23755.500011574073, 23755.50695601852, 23755.513900462964, 23755.52084490741, 23755.52778935185, 23755.534733796296, 23755.54167824074, 23755.548622685186, 23755.555567129628, 23755.562511574073, 23755.56945601852, 23755.576400462964, 23755.58334490741, 23755.59028935185, 23755.597233796296, 23755.60417824074, 23755.611122685186, 23755.618067129628, 23755.625011574073, 23755.63195601852, 23755.638900462964, 23755.64584490741, 23755.65278935185, 23755.659733796296, 23755.66667824074, 23755.673622685186, 23755.680567129628, 23755.687511574073, 23755.69445601852, 23755.701400462964, 23755.70834490741, 23755.71528935185, 23755.722233796296, 23755.72917824074, 23755.736122685186, 23755.743067129628, 23755.750011574073, 23755.75695601852, 23755.763900462964, 23755.77084490741, 23755.77778935185, 23755.784733796296, 23755.79167824074, 23755.798622685186, 23755.805567129628, 23755.812511574073, 23755.81945601852, 23755.826400462964, 23755.83334490741, 23755.84028935185, 23755.847233796296, 23755.85417824074, 23755.861122685186, 23755.868067129628, 23755.875011574073, 23755.88195601852, 23755.888900462964, 23755.89584490741, 23755.90278935185, 23755.909733796296, 23755.91667824074, 23755.923622685186, 23755.930567129628, 23755.937511574073, 23755.94445601852, 23755.951400462964, 23755.95834490741, 23755.96528935185, 23755.972233796296, 23755.97917824074, 23755.986122685186, 23755.993067129628, 23756.000011574073, 23756.00695601852, 23756.013900462964, 23756.02084490741, 23756.02778935185, 23756.034733796296, 23756.04167824074, 23756.048622685186, 23756.055567129628, 23756.062511574073, 23756.06945601852, 23756.076400462964, 23756.08334490741, 23756.09028935185, 23756.097233796296, 23756.10417824074, 23756.111122685186, 23756.118067129628, 23756.125011574073, 23756.13195601852, 23756.138900462964, 23756.14584490741, 23756.15278935185, 23756.159733796296, 23756.16667824074, 23756.173622685186, 23756.180567129628, 23756.187511574073, 23756.19445601852, 23756.201400462964, 23756.20834490741, 23756.21528935185, 23756.222233796296, 23756.22917824074, 23756.236122685186, 23756.243067129628, 23756.250011574073, 23756.25695601852, 23756.263900462964, 23756.27084490741, 23756.27778935185, 23756.284733796296, 23756.29167824074, 23756.298622685186, 23756.305567129628, 23756.312511574073, 23756.31945601852, 23756.326400462964, 23756.33334490741, 23756.34028935185, 23756.347233796296, 23756.35417824074, 23756.361122685186, 23756.368067129628, 23756.375011574073, 23756.38195601852, 23756.388900462964, 23756.39584490741, 23756.40278935185, 23756.409733796296, 23756.41667824074, 23756.423622685186, 23756.430567129628, 23756.437511574073, 23756.44445601852, 23756.451400462964, 23756.45834490741, 23756.46528935185, 23756.472233796296, 23756.47917824074, 23756.486122685186, 23756.493067129628, 23756.500011574073, 23756.50695601852, 23756.513900462964, 23756.52084490741, 23756.52778935185, 23756.534733796296, 23756.54167824074, 23756.548622685186, 23756.555567129628, 23756.562511574073, 23756.56945601852, 23756.576400462964, 23756.58334490741, 23756.59028935185, 23756.597233796296, 23756.60417824074, 23756.611122685186, 23756.618067129628, 23756.625011574073, 23756.63195601852, 23756.638900462964, 23756.64584490741, 23756.65278935185, 23756.659733796296, 23756.66667824074, 23756.673622685186, 23756.680567129628, 23756.687511574073, 23756.69445601852, 23756.701400462964, 23756.70834490741, 23756.71528935185, 23756.722233796296, 23756.72917824074, 23756.736122685186, 23756.743067129628, 23756.750011574073, 23756.75695601852, 23756.763900462964, 23756.77084490741, 23756.77778935185, 23756.784733796296, 23756.79167824074, 23756.798622685186, 23756.805567129628, 23756.812511574073, 23756.81945601852, 23756.826400462964, 23756.83334490741, 23756.84028935185, 23756.847233796296, 23756.85417824074, 23756.861122685186, 23756.868067129628, 23756.875011574073, 23756.88195601852, 23756.888900462964, 23756.89584490741, 23756.90278935185, 23756.909733796296, 23756.91667824074, 23756.923622685186, 23756.930567129628, 23756.937511574073, 23756.94445601852, 23756.951400462964, 23756.95834490741, 23756.96528935185, 23756.972233796296, 23756.97917824074, 23756.986122685186, 23756.993067129628, 23757.000011574073, 23757.00695601852, 23757.013900462964, 23757.02084490741, 23757.02778935185, 23757.034733796296, 23757.04167824074, 23757.048622685186, 23757.055567129628, 23757.062511574073, 23757.06945601852, 23757.076400462964, 23757.08334490741, 23757.09028935185, 23757.097233796296, 23757.10417824074, 23757.111122685186, 23757.118067129628, 23757.125011574073, 23757.13195601852, 23757.138900462964, 23757.14584490741, 23757.15278935185, 23757.159733796296, 23757.16667824074, 23757.173622685186, 23757.180567129628, 23757.187511574073, 23757.19445601852, 23757.201400462964, 23757.20834490741, 23757.21528935185, 23757.222233796296, 23757.22917824074, 23757.236122685186, 23757.243067129628, 23757.250011574073, 23757.25695601852, 23757.263900462964, 23757.27084490741, 23757.27778935185, 23757.284733796296, 23757.29167824074, 23757.298622685186, 23757.305567129628, 23757.312511574073, 23757.31945601852, 23757.326400462964, 23757.33334490741, 23757.34028935185, 23757.347233796296, 23757.35417824074, 23757.361122685186, 23757.368067129628, 23757.375011574073, 23757.38195601852, 23757.388900462964, 23757.39584490741, 23757.40278935185, 23757.409733796296, 23757.41667824074, 23757.423622685186, 23757.430567129628, 23757.437511574073, 23757.44445601852, 23757.451400462964, 23757.45834490741, 23757.46528935185, 23757.472233796296, 23757.47917824074, 23757.486122685186, 23757.493067129628, 23757.500011574073, 23757.50695601852, 23757.513900462964, 23757.52084490741, 23757.52778935185, 23757.534733796296, 23757.54167824074, 23757.548622685186, 23757.555567129628, 23757.562511574073, 23757.56945601852, 23757.576400462964, 23757.58334490741, 23757.59028935185, 23757.597233796296, 23757.60417824074, 23757.611122685186, 23757.618067129628, 23757.625011574073, 23757.63195601852, 23757.638900462964, 23757.64584490741, 23757.65278935185, 23757.659733796296, 23757.66667824074, 23757.673622685186, 23757.680567129628, 23757.687511574073, 23757.69445601852, 23757.701400462964, 23757.70834490741, 23757.71528935185, 23757.722233796296, 23757.72917824074, 23757.736122685186, 23757.743067129628, 23757.750011574073, 23757.75695601852, 23757.763900462964, 23757.77084490741, 23757.77778935185, 23757.784733796296, 23757.79167824074, 23757.798622685186, 23757.805567129628, 23757.812511574073, 23757.81945601852, 23757.826400462964, 23757.83334490741, 23757.84028935185, 23757.847233796296, 23757.85417824074, 23757.861122685186, 23757.868067129628, 23757.875011574073, 23757.88195601852, 23757.888900462964, 23757.89584490741, 23757.90278935185, 23757.909733796296, 23757.91667824074, 23757.923622685186, 23757.930567129628, 23757.937511574073, 23757.94445601852, 23757.951400462964, 23757.95834490741, 23757.96528935185, 23757.972233796296, 23757.97917824074, 23757.986122685186, 23757.993067129628, 23758.000011574073, 23758.00695601852, 23758.013900462964, 23758.02084490741, 23758.02778935185, 23758.034733796296, 23758.04167824074, 23758.048622685186, 23758.055567129628, 23758.062511574073, 23758.06945601852, 23758.076400462964, 23758.08334490741, 23758.09028935185, 23758.097233796296, 23758.10417824074, 23758.111122685186, 23758.118067129628, 23758.125011574073, 23758.13195601852, 23758.138900462964, 23758.14584490741, 23758.15278935185, 23758.159733796296, 23758.16667824074, 23758.173622685186, 23758.180567129628, 23758.187511574073, 23758.19445601852, 23758.201400462964, 23758.20834490741, 23758.21528935185, 23758.222233796296, 23758.22917824074, 23758.236122685186, 23758.243067129628, 23758.250011574073, 23758.25695601852, 23758.263900462964, 23758.27084490741, 23758.27778935185, 23758.284733796296, 23758.29167824074, 23758.298622685186, 23758.305567129628, 23758.312511574073, 23758.31945601852, 23758.326400462964, 23758.33334490741, 23758.34028935185, 23758.347233796296, 23758.35417824074, 23758.361122685186, 23758.368067129628, 23758.375011574073, 23758.38195601852, 23758.388900462964, 23758.39584490741, 23758.40278935185, 23758.409733796296, 23758.41667824074, 23758.423622685186, 23758.430567129628, 23758.437511574073, 23758.44445601852, 23758.451400462964, 23758.45834490741, 23758.46528935185, 23758.472233796296, 23758.47917824074, 23758.486122685186, 23758.493067129628, 23758.500011574073, 23758.50695601852, 23758.513900462964, 23758.52084490741, 23758.52778935185, 23758.534733796296, 23758.54167824074, 23758.548622685186, 23758.555567129628, 23758.562511574073, 23758.56945601852, 23758.576400462964, 23758.58334490741, 23758.59028935185, 23758.597233796296, 23758.60417824074, 23758.611122685186, 23758.618067129628, 23758.625011574073, 23758.63195601852, 23758.638900462964, 23758.64584490741, 23758.65278935185, 23758.659733796296, 23758.66667824074, 23758.673622685186, 23758.680567129628, 23758.687511574073, 23758.69445601852, 23758.701400462964, 23758.70834490741, 23758.71528935185, 23758.722233796296, 23758.72917824074, 23758.736122685186, 23758.743067129628, 23758.750011574073, 23758.75695601852, 23758.763900462964, 23758.77084490741, 23758.77778935185, 23758.784733796296, 23758.79167824074, 23758.798622685186, 23758.805567129628, 23758.812511574073, 23758.81945601852, 23758.826400462964, 23758.83334490741, 23758.84028935185, 23758.847233796296, 23758.85417824074, 23758.861122685186, 23758.868067129628, 23758.875011574073, 23758.88195601852, 23758.888900462964, 23758.89584490741, 23758.90278935185, 23758.909733796296, 23758.91667824074, 23758.923622685186, 23758.930567129628, 23758.937511574073, 23758.94445601852, 23758.951400462964, 23758.95834490741, 23758.96528935185, 23758.972233796296, 23758.97917824074, 23758.986122685186, 23758.993067129628, 23759.000011574073, 23759.00695601852, 23759.013900462964, 23759.02084490741, 23759.02778935185, 23759.034733796296, 23759.04167824074, 23759.048622685186, 23759.055567129628, 23759.062511574073, 23759.06945601852, 23759.076400462964, 23759.08334490741, 23759.09028935185, 23759.097233796296, 23759.10417824074, 23759.111122685186, 23759.118067129628, 23759.125011574073, 23759.13195601852, 23759.138900462964, 23759.14584490741, 23759.15278935185, 23759.159733796296, 23759.16667824074, 23759.173622685186, 23759.180567129628, 23759.187511574073, 23759.19445601852, 23759.201400462964, 23759.20834490741, 23759.21528935185, 23759.222233796296, 23759.22917824074, 23759.236122685186, 23759.243067129628, 23759.250011574073, 23759.25695601852, 23759.263900462964, 23759.27084490741, 23759.27778935185, 23759.284733796296, 23759.29167824074, 23759.298622685186, 23759.305567129628, 23759.312511574073, 23759.31945601852, 23759.326400462964, 23759.33334490741, 23759.34028935185, 23759.347233796296, 23759.35417824074, 23759.361122685186, 23759.368067129628, 23759.375011574073, 23759.38195601852, 23759.388900462964, 23759.39584490741, 23759.40278935185, 23759.409733796296, 23759.41667824074, 23759.423622685186, 23759.430567129628, 23759.437511574073, 23759.44445601852, 23759.451400462964, 23759.45834490741, 23759.46528935185, 23759.472233796296, 23759.47917824074, 23759.486122685186, 23759.493067129628, 23759.500011574073, 23759.50695601852, 23759.513900462964, 23759.52084490741, 23759.52778935185, 23759.534733796296, 23759.54167824074, 23759.548622685186, 23759.555567129628, 23759.562511574073, 23759.56945601852, 23759.576400462964, 23759.58334490741, 23759.59028935185, 23759.597233796296, 23759.60417824074, 23759.611122685186, 23759.618067129628, 23759.625011574073, 23759.63195601852, 23759.638900462964, 23759.64584490741, 23759.65278935185, 23759.659733796296, 23759.66667824074, 23759.673622685186, 23759.680567129628, 23759.687511574073, 23759.69445601852, 23759.701400462964, 23759.70834490741, 23759.71528935185, 23759.722233796296, 23759.72917824074, 23759.736122685186, 23759.743067129628, 23759.750011574073, 23759.75695601852, 23759.763900462964, 23759.77084490741, 23759.77778935185, 23759.784733796296, 23759.79167824074, 23759.798622685186, 23759.805567129628, 23759.812511574073, 23759.81945601852, 23759.826400462964, 23759.83334490741, 23759.84028935185, 23759.847233796296, 23759.85417824074, 23759.861122685186, 23759.868067129628, 23759.875011574073, 23759.88195601852, 23759.888900462964, 23759.89584490741, 23759.90278935185, 23759.909733796296, 23759.91667824074, 23759.923622685186, 23759.930567129628, 23759.937511574073, 23759.94445601852, 23759.951400462964, 23759.95834490741, 23759.96528935185, 23759.972233796296, 23759.97917824074, 23759.986122685186, 23759.993067129628, 23760.000011574073, 23760.00695601852, 23760.013900462964, 23760.02084490741, 23760.02778935185, 23760.034733796296, 23760.04167824074, 23760.048622685186, 23760.055567129628, 23760.062511574073, 23760.06945601852, 23760.076400462964, 23760.08334490741, 23760.09028935185, 23760.097233796296, 23760.10417824074, 23760.111122685186, 23760.118067129628, 23760.125011574073, 23760.13195601852, 23760.138900462964, 23760.14584490741, 23760.15278935185, 23760.159733796296, 23760.16667824074, 23760.173622685186, 23760.180567129628, 23760.187511574073, 23760.19445601852, 23760.201400462964, 23760.20834490741, 23760.21528935185, 23760.222233796296, 23760.22917824074, 23760.236122685186, 23760.243067129628, 23760.250011574073, 23760.25695601852, 23760.263900462964, 23760.27084490741, 23760.27778935185, 23760.284733796296, 23760.29167824074, 23760.298622685186, 23760.305567129628, 23760.312511574073, 23760.31945601852, 23760.326400462964, 23760.33334490741, 23760.34028935185, 23760.347233796296, 23760.35417824074, 23760.361122685186, 23760.368067129628, 23760.375011574073, 23760.38195601852, 23760.388900462964, 23760.39584490741, 23760.40278935185, 23760.409733796296, 23760.41667824074, 23760.423622685186, 23760.430567129628, 23760.437511574073, 23760.44445601852, 23760.451400462964, 23760.45834490741, 23760.46528935185, 23760.472233796296, 23760.47917824074, 23760.486122685186, 23760.493067129628, 23760.500011574073, 23760.50695601852, 23760.513900462964, 23760.52084490741, 23760.52778935185, 23760.534733796296, 23760.54167824074, 23760.548622685186, 23760.555567129628, 23760.562511574073, 23760.56945601852, 23760.576400462964, 23760.58334490741, 23760.59028935185, 23760.597233796296, 23760.60417824074, 23760.611122685186, 23760.618067129628, 23760.625011574073, 23760.63195601852, 23760.638900462964, 23760.64584490741, 23760.65278935185, 23760.659733796296, 23760.66667824074, 23760.673622685186, 23760.680567129628, 23760.687511574073, 23760.69445601852, 23760.701400462964, 23760.70834490741, 23760.71528935185, 23760.722233796296, 23760.72917824074, 23760.736122685186, 23760.743067129628, 23760.750011574073, 23760.75695601852, 23760.763900462964, 23760.77084490741, 23760.77778935185, 23760.784733796296, 23760.79167824074, 23760.798622685186, 23760.805567129628, 23760.812511574073, 23760.81945601852, 23760.826400462964, 23760.83334490741, 23760.84028935185, 23760.847233796296, 23760.85417824074, 23760.861122685186, 23760.868067129628, 23760.875011574073, 23760.88195601852, 23760.888900462964, 23760.89584490741, 23760.90278935185, 23760.909733796296, 23760.91667824074, 23760.923622685186, 23760.930567129628, 23760.937511574073, 23760.94445601852, 23760.951400462964, 23760.95834490741, 23760.96528935185, 23760.972233796296, 23760.97917824074, 23760.986122685186, 23760.993067129628, 23761.000011574073, 23761.00695601852, 23761.013900462964, 23761.02084490741, 23761.02778935185, 23761.034733796296, 23761.04167824074, 23761.048622685186, 23761.055567129628, 23761.062511574073, 23761.06945601852, 23761.076400462964, 23761.08334490741, 23761.09028935185, 23761.097233796296, 23761.10417824074, 23761.111122685186, 23761.118067129628, 23761.125011574073, 23761.13195601852, 23761.138900462964, 23761.14584490741, 23761.15278935185, 23761.159733796296, 23761.16667824074, 23761.173622685186, 23761.180567129628, 23761.187511574073, 23761.19445601852, 23761.201400462964, 23761.20834490741}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =70.0
TEMP =
  {19.6662, 19.6179, 19.5821, 19.6573, 19.7039, 19.6881, 19.7673, 19.7747, 19.7157, 19.6752, 19.7103, 19.7358, 19.6427, 19.6064, 19.5894, 19.659, 19.6879, 19.6966, 19.7321, 19.7888, 19.7907, 19.8199, 19.8597, 19.8818, 19.9025, 19.9276, 19.9339, 19.7923, 19.9124, 19.8328, 19.8442, 19.7283, 19.6258, 19.6595, 19.7141, 19.8578, 19.8791, 19.7657, 19.7038, 19.5779, 19.6937, 19.7018, 19.668, 19.6993, 19.8086, 19.6564, 19.6861, 19.6641, 19.6855, 19.6958, 19.7697, 19.7296, 19.6687, 19.663, 19.5356, 19.5754, 19.5392, 19.4632, 19.5103, 19.398, 19.3789, 19.4719, 19.6637, 19.6861, 19.6031, 19.5414, 19.512, 19.4487, 19.4479, 19.4621, 19.4577, 19.491, 19.5656, 19.7428, 19.742, 19.7753, 19.7673, 19.7204, 19.754, 19.7604, 19.932, 19.8727, 19.9719, 19.9102, 19.9041, 19.8562, 19.9618, 19.9411, 19.8897, 19.8924, 19.8925, 20.079, 20.1487, 20.1324, 20.1353, 20.1092, 20.0098, 19.8966, 19.9063, 19.743, 19.7295, 19.7655, 19.7653, 19.6984, 19.6856, 19.6725, 19.6692, 19.6397, 19.6896, 19.5693, 19.5655, 19.5395, 19.5774, 19.464, 19.62, 19.6019, 19.6089, 19.6567, 19.6352, 19.6296, 19.6216, 19.5955, 19.6253, 19.6548, 19.5791, 19.6844, 19.602, 19.5942, 19.6051, 19.5639, 19.5961, 19.6241, 19.6161, 19.5571, 19.5303, 19.5276, 19.5433, 19.5367, 19.5112, 19.5411, 19.5051, 19.5183, 19.4901, 19.4554, 19.4783, 19.5454, 19.5487, 19.5886, 19.5942, 19.6045, 19.6718, 19.6729, 19.6614, 19.7438, 19.7818, 19.7711, 19.6847, 19.8453, 19.698, 19.7024, 19.6893, 19.7026, 19.8978, 19.8775, 19.7432, 19.6457, 19.6127, 19.2728, 19.3471, 19.4154, 19.2322, 19.0823, 19.3694, 19.6641, 19.4354, 19.6745, 19.4741, 19.4579, 19.0522, 19.015, 19.7453, 19.7642, 19.711, 19.9063, 19.8536, 19.0417, 18.9663, 18.9465, 18.946, 18.9558, 18.9737, 18.963, 18.9538, 18.9519, 18.9581, 18.977, 18.972, 18.9788, 18.9824, 19.1012, 19.1718, 19.017, 18.9537, 18.9882, 19.0017, 19.0047, 18.9437, 18.8947, 18.8768, 18.9223, 18.9878, 18.9819, 18.9453, 19.08, 19.2026, 19.0559, 19.0861, 19.1361, 19.2086, 19.2515, 19.2164, 19.2312, 19.2236, 19.2786, 19.3243, 19.3204, 19.3295, 19.396, 19.4124, 19.4669, 19.4565, 19.6275, 19.894, 19.4614, 19.4575, 19.4629, 19.5036, 19.5118, 19.4704, 19.4579, 19.5127, 19.4933, 19.4369, 19.3512, 19.3471, 19.3649, 19.343, 19.1772, 19.1791, 19.2925, 19.3309, 19.3431, 19.312, 19.1739, 19.1221, 18.9338, 19.131, 19.1003, 19.1508, 19.1401, 19.1369, 19.2536, 19.3486, 19.2579, 19.1448, 18.9586, 18.9468, 18.9465, 18.9652, 18.9698, 18.8872, 18.8195, 18.9769, 19.2827, 19.2298, 19.3234, 19.2447, 19.3134, 18.929, 18.8655, 19.226, 19.2739, 19.0702, 18.8608, 18.8302, 18.8925, 18.9645, 19.0735, 18.9032, 19.0227, 18.9653, 18.7657, 18.7239, 18.7519, 18.5123, 18.4417, 18.505, 18.4646, 18.4266, 18.3052, 18.2949, 18.2874, 18.2919, 18.5638, 18.7662, 18.787, 18.7529, 18.7363, 18.7776, 18.7667, 18.7591, 18.8769, 18.775, 18.7726, 18.7757, 18.7891, 18.7958, 18.9459, 18.8684, 18.8028, 18.8175, 18.9148, 19.2474, 19.1814, 19.1536, 19.0071, 18.889, 19.1616, 19.0917, 18.9983, 19.1366, 19.0822, 19.1209, 19.3298, 19.3018, 18.993, 18.993, 18.9552, 18.9572, 19.155, 19.1797, 19.1465, 19.1494, 19.1881, 19.1046, 18.9805, 18.925, 18.9345, 18.8757, 19.3112, 19.1598, 19.0392, 19.0228, 19.0109, 18.8257, 18.8285, 18.8381, 19.0317, 18.9327, 19.0371, 18.8079, 19.1488, 19.237, 18.8275, 19.1538, 18.9355, 19.0503, 19.2009, 19.3787, 19.0588, 19.1967, 19.1639, 19.2465, 19.2584, 19.1557, 18.9724, 19.199, 19.3732, 19.4295, 19.2832, 19.4237, 19.4541, 19.419, 19.4515, 19.4116, 19.3658, 19.4572, 19.3713, 19.3887, 19.1126, 19.0325, 19.2441, 19.083, 19.1508, 19.0064, 18.9877, 19.0745, 19.026, 19.0094, 19.169, 19.2248, 19.3549, 19.3208, 19.3248, 19.2812, 19.3052, 19.2829, 19.3286, 19.3631, 19.3994, 19.2994, 19.2243, 18.9717, 18.8031, 19.0919, 19.205, 19.4158, 19.1024, 18.8161, 18.8327, 18.8086, 18.8045, 18.7667, 18.7291, 18.6146, 18.487, 18.5149, 18.5491, 18.9044, 18.8992, 18.9087, 18.8213, 18.5594, 18.9587, 18.7846, 18.8935, 18.8474, 18.8187, 18.6182, 18.5485, 18.5003, 18.476, 18.4024, 18.501, 18.515, 18.54, 18.5518, 18.5461, 18.5286, 18.533, 18.5462, 18.6708, 18.6609, 18.5944, 18.5454, 18.569, 18.6023, 18.5921, 18.5904, 18.6202, 18.6324, 18.6191, 18.6227, 18.6361, 18.6269, 18.6234, 18.6472, 18.6521, 18.6609, 18.6765, 18.7293, 18.6925, 18.7599, 18.8335, 18.8108, 18.8951, 18.8312, 18.9146, 19.0451, 19.1373, 19.1222, 18.9738, 19.1615, 19.1805, 19.0959, 18.7829, 18.8383, 19.0244, 18.9371, 18.9217, 18.9024, 18.8965, 18.8484, 18.8351, 18.9131, 18.9854, 18.8825, 18.9096, 18.9225, 19.014, 18.9516, 18.9718, 19.2411, 19.2988, 19.319, 19.2948, 19.4473, 19.4482, 19.6192, 19.5352, 19.6172, 19.5937, 19.4516, 19.3382, 19.1144, 19.1525, 19.1804, 19.3244, 19.241, 19.2209, 19.1686, 19.2372, 19.2369, 19.5341, 19.5222, 19.5416, 19.4366, 19.5447, 19.5786, 19.7105, 19.6859, 19.2957, 19.284, 19.3059, 19.6031, 19.3183, 19.3065, 19.3171, 19.3294, 19.2638, 19.2628, 19.2756, 19.3052, 19.5623, 19.5506, 19.5671, 19.5914, 19.5877, 19.6019, 19.6641, 19.3995, 19.3921, 19.3603, 19.6243, 19.706, 19.3378, 19.1971, 19.1938, 19.2703, 19.2602, 19.379, 19.3405, 19.2156, 19.1716, 19.2586, 19.2394, 19.2424, 19.1695, 18.9897, 19.1865, 19.2209, 19.3155, 19.3366, 19.0148, 18.9278, 18.965, 18.8583, 18.9148, 19.0846, 19.0832, 18.8929, 18.8244, 18.7532, 18.729, 18.5837, 18.5884, 18.6114, 18.8206, 18.9373, 18.9999, 18.7103, 18.8087, 18.7709, 18.7049, 18.6887, 18.7395, 18.9153, 18.8279, 18.776, 18.7534, 18.8859, 19.1089, 19.0359, 19.165, 19.0195, 18.7973, 18.7199, 18.707, 18.6318, 18.6015, 18.6591, 18.6583, 18.6426, 18.663, 18.6569, 18.5251, 18.4569, 18.466, 18.5424, 18.5896, 18.4978, 18.4792, 18.4607, 18.4548, 18.4321, 18.4323, 18.4255, 18.4223, 18.4216, 18.4308, 18.4408, 18.4398, 18.4352, 18.4607, 18.4648, 18.4709, 18.4689, 18.4763, 18.4909, 18.5002, 18.4811, 18.5028, 18.5154, 18.6612, 18.556, 18.5799, 18.8166, 18.7938, 18.9512, 18.7855, 18.8507, 18.9386, 18.9155, 18.8489, 18.7434, 18.7287, 18.7087, 18.7529, 18.7325, 18.7515, 18.7794, 18.8171, 18.8128, 18.8301, 18.9486, 19.0552, 19.23, 19.4404, 19.4073, 19.3308, 19.392, 19.0463, 19.0815, 19.1014, 19.0763, 18.9598, 18.9313, 18.9691, 18.997, 19.0146, 19.0796, 19.1069, 19.0451, 19.0306, 18.9656, 19.0953, 19.1366, 19.1232, 18.9789, 18.9256, 19.0316, 18.9063, 19.0481, 19.2512, 19.0337, 18.9501, 18.8781, 18.8279, 18.8799, 18.8455, 18.8057, 18.8069, 18.8067, 18.8126, 18.7266, 18.7984, 18.8828, 19.0601, 19.048, 19.1533, 19.4497, 19.2888, 19.3258, 19.2308, 19.0294, 18.9455, 18.8929, 18.9083, 18.9405, 19.2589, 19.0804, 18.996, 18.8975, 18.8469, 18.5815, 18.9399, 18.8677, 18.5575, 18.5079, 18.6184, 18.5894, 18.6415, 18.6401, 18.6671, 18.5922, 18.6133, 18.5722, 18.5179, 18.5327, 18.6149, 18.5684, 18.752, 18.6294, 18.6406, 18.6365, 18.7411, 18.7189, 18.8852, 18.9016, 18.8939, 18.9055, 18.9107, 18.8124, 18.8071, 18.7673, 18.8876, 18.926, 18.8914, 18.8208, 18.7041, 18.685, 18.6371, 18.6799, 18.7192, 18.6915, 18.7078, 18.6963, 18.7856, 18.7779, 18.7813, 18.7705, 18.787, 18.7673, 18.7935, 18.667, 18.7353, 18.7627, 18.7708, 18.7907, 18.7669, 18.7959, 18.8154, 18.8064, 18.783, 18.7946, 18.811, 18.8119, 18.8103, 18.8079, 19.4362, 18.8296, 19.4449, 19.0144, 19.2269, 19.254, 18.8492, 18.7096, 18.9878, 18.6815, 18.8364, 18.6419, 18.6807, 18.9691, 18.8964, 19.3236, 18.9475, 18.9078, 18.957, 18.7701, 18.7817, 18.6957, 18.8997, 18.8235, 18.8805, 19.2089, 19.3637, 19.6882, 18.8721, 19.1008, 18.8004, 19.0489, 18.8432, 18.9005, 18.8502, 18.7529, 18.743, 18.9097, 18.9706, 19.2918, 18.9913, 18.9575, 19.2064, 19.2462, 19.278, 19.1014, 19.0683, 19.017, 18.9634, 19.0771, 19.0158, 19.0674, 18.9649, 18.7994, 18.8105, 19.0194, 19.0214, 18.8247, 18.8167, 19.1249, 18.9037, 18.9587, 18.9262, 18.8271, 18.8006, 18.7901, 18.7698, 18.768, 18.7599, 18.909, 18.9162, 18.9451, 18.8526, 18.8247, 18.6358, 18.7552, 18.8028, 18.7475, 18.8225, 18.8049, 18.5764, 18.5845, 18.5008, 18.4454, 18.6739, 18.4612, 18.4497, 18.4329, 18.3174, 18.2818, 18.3272, 18.3809, 18.416, 18.3706, 18.4363, 18.368, 18.4444, 18.4947, 22.6714, 24.9047, 22.4275, 24.0492, 22.8552, 22.8845, 24.41, 22.2899, 22.1926, 21.9761, 21.7615, 21.7765, 21.7783, 21.7748, 21.9514, 22.1062, 22.5306, 23.3426, 23.8617, 23.375, 27.3326, 27.9231, 27.8623, 27.8226, 27.7966, 27.758, 27.7081, 27.6643, 27.6154, 27.5667, 27.5112, 27.4483, 27.3812, 27.3146, 27.2372, 27.1641, 27.0931, 27.0215, 26.9436, 26.8721, 26.7979, 26.7247, 26.6573, 26.5886, 26.5174, 26.4446, 26.375, 26.3061, 26.2387, 26.1584, 26.0946, 26.0248, 25.9498, 25.8679, 25.787, 25.7145, 25.6254, 25.5447, 25.4757, 25.3993, 25.329, 25.2563, 25.1831, 25.1169, 25.0472, 24.9785, 24.9168, 24.8466, 24.7886, 24.7336, 24.6683, 24.6131, 24.561, 24.499, 24.4397, 24.3845, 24.328, 24.2564, 24.1903, 24.1165, 24.0452, 23.967, 23.8927, 23.8229, 23.7607, 23.6968, 23.6468, 23.5985, 23.5555, 23.5119, 23.4619, 23.4168, 23.3705, 23.3093, 23.2558, 23.1968, 23.1456, 23.0812, 23.0304, 22.976, 22.9161, 22.8556, 22.7916, 22.7414, 22.6865, 22.6203, 22.571, 22.5095, 22.458, 22.408, 22.3492, 22.2903, 22.2381, 22.175, 22.1206, 22.0713, 22.017, 21.9616, 21.9121, 21.8621, 21.8152, 21.7692, 21.7299, 21.6909, 21.6427, 21.6107, 21.5684, 21.5393, 21.5044, 21.4747, 21.4467, 21.4195, 21.3961, 21.3779, 21.3637, 21.3528, 21.3447, 21.3395, 21.3368, 21.3363, 21.3391, 21.3472, 21.3545, 21.3697, 21.3826, 21.3923, 21.4066, 21.4265, 21.441, 21.4744, 24.1563, 23.4123, 23.4489, 23.443, 23.2704, 23.3133, 23.6231, 23.7617}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {4.848557, 4.8439536, 4.8399963, 4.847583, 4.852098, 4.850581, 4.8581467, 4.8588543, 4.8534985, 4.849497, 4.8527503, 4.8554277, 4.8475485, 4.844139, 4.8421154, 4.849051, 4.8517485, 4.852778, 4.8561764, 4.8614507, 4.862021, 4.8645773, 4.868027, 4.87, 4.8721037, 4.874621, 4.8753843, 4.863395, 4.874779, 4.866556, 4.8674774, 4.8565335, 4.846554, 4.8491197, 4.8546314, 4.870626, 4.8732595, 4.861135, 4.8542953, 4.8411627, 4.8539176, 4.8552637, 4.851529, 4.855181, 4.8662543, 4.8509593, 4.8536844, 4.851783, 4.8538423, 4.854879, 4.862578, 4.8585596, 4.852188, 4.851282, 4.8384614, 4.841327, 4.837522, 4.8284693, 4.8340607, 4.8217316, 4.8199105, 4.8289285, 4.848365, 4.851007, 4.8422937, 4.83587, 4.8327923, 4.826579, 4.8265724, 4.8281546, 4.8280654, 4.8313055, 4.8380017, 4.8562245, 4.856094, 4.8602695, 4.859775, 4.8545904, 4.858573, 4.860297, 4.882169, 4.874807, 4.887001, 4.8805037, 4.880579, 4.87608, 4.8866706, 4.8848395, 4.879616, 4.8801045, 4.8799186, 4.898705, 4.9064474, 4.904565, 4.9049025, 4.9022064, 4.8914843, 4.878164, 4.879946, 4.8616576, 4.8590884, 4.862743, 4.8628187, 4.855984, 4.854735, 4.8533344, 4.852957, 4.849978, 4.8545904, 4.842932, 4.842514, 4.8396406, 4.8433986, 4.8327107, 4.847432, 4.8461423, 4.846835, 4.8517075, 4.849745, 4.849072, 4.8482623, 4.845731, 4.848777, 4.852154, 4.8452096, 4.855325, 4.8480635, 4.8477616, 4.848997, 4.845539, 4.8484893, 4.8514333, 4.85061, 4.843817, 4.840772, 4.8403673, 4.8417597, 4.840765, 4.8380294, 4.8409367, 4.837337, 4.838331, 4.8356028, 4.8325877, 4.834294, 4.841197, 4.841581, 4.8452644, 4.8458953, 4.847137, 4.85365, 4.8541307, 4.8527784, 4.860737, 4.864756, 4.8638215, 4.855044, 4.871059, 4.856616, 4.856561, 4.8547964, 4.856204, 4.8760724, 4.8748345, 4.860579, 4.850616, 4.8477545, 4.814081, 4.819815, 4.82571, 4.8083563, 4.7942867, 4.82128, 4.850616, 4.8297167, 4.853046, 4.8318677, 4.830258, 4.7917876, 4.787043, 4.858903, 4.863671, 4.856218, 4.876719, 4.871623, 4.7924366, 4.782192, 4.779798, 4.779661, 4.7807393, 4.7826014, 4.781585, 4.780603, 4.7803845, 4.780971, 4.782956, 4.7825127, 4.783195, 4.7835975, 4.795837, 4.803107, 4.7871118, 4.7806234, 4.784109, 4.785638, 4.78589, 4.779757, 4.774288, 4.7726116, 4.777268, 4.78428, 4.783727, 4.7799206, 4.792996, 4.805478, 4.791822, 4.7943687, 4.7992387, 4.8059907, 4.8104625, 4.8072968, 4.8084316, 4.8077, 4.8132257, 4.817276, 4.817016, 4.817885, 4.824395, 4.826532, 4.8321967, 4.8319845, 4.848269, 4.8768086, 4.8320665, 4.830881, 4.8313265, 4.835651, 4.836439, 4.8322515, 4.8310733, 4.8363976, 4.8349037, 4.829689, 4.821424, 4.820986, 4.822594, 4.820609, 4.8039675, 4.8042684, 4.816099, 4.819398, 4.8202395, 4.817666, 4.803407, 4.798091, 4.778802, 4.79889, 4.795789, 4.8007145, 4.7999153, 4.7994165, 4.810996, 4.8201094, 4.811796, 4.800496, 4.780964, 4.779327, 4.779238, 4.7816596, 4.7816734, 4.773211, 4.7663765, 4.781987, 4.813397, 4.8089857, 4.8176866, 4.8105516, 4.8170915, 4.779034, 4.771146, 4.8076863, 4.813274, 4.7930846, 4.7708187, 4.767528, 4.77362, 4.780732, 4.7932487, 4.7748747, 4.7883744, 4.7810526, 4.7611327, 4.7561154, 4.7593894, 4.7353697, 4.7271867, 4.733536, 4.7295017, 4.725999, 4.713266, 4.7123914, 4.711449, 4.711815, 4.7392154, 4.7607036, 4.7628894, 4.7594576, 4.7571363, 4.761936, 4.760867, 4.760118, 4.7718344, 4.7618613, 4.7614865, 4.762147, 4.763169, 4.7638974, 4.779034, 4.7715144, 4.7647963, 4.766138, 4.7758837, 4.809895, 4.803913, 4.8005643, 4.786061, 4.7739134, 4.801405, 4.794075, 4.7849073, 4.798904, 4.793351, 4.7975583, 4.8183026, 4.8157983, 4.784628, 4.784075, 4.780439, 4.7804866, 4.800086, 4.803086, 4.7996078, 4.799936, 4.803236, 4.7955227, 4.78355, 4.777138, 4.7779837, 4.7728233, 4.815518, 4.8015757, 4.7889066, 4.78761, 4.786675, 4.7671876, 4.767644, 4.76823, 4.788811, 4.7784133, 4.789303, 4.7653823, 4.8003116, 4.809649, 4.7680936, 4.801583, 4.7789044, 4.790791, 4.806285, 4.8249774, 4.791849, 4.806121, 4.8028607, 4.810538, 4.8132057, 4.801528, 4.782717, 4.806169, 4.824498, 4.8308268, 4.815463, 4.829799, 4.8333344, 4.829696, 4.8329577, 4.8288813, 4.8237314, 4.8334236, 4.824313, 4.826614, 4.7980366, 4.789371, 4.8105173, 4.794341, 4.8013363, 4.786327, 4.784198, 4.792914, 4.7885246, 4.7865863, 4.802703, 4.808452, 4.821944, 4.818515, 4.8189735, 4.814245, 4.8167424, 4.814457, 4.819131, 4.8227863, 4.8267236, 4.816236, 4.807871, 4.7826214, 4.7656, 4.793986, 4.806394, 4.828751, 4.797285, 4.766438, 4.7678347, 4.765205, 4.765116, 4.7613845, 4.757375, 4.74553, 4.7323337, 4.734867, 4.7386446, 4.775236, 4.775004, 4.7761016, 4.7663083, 4.7401056, 4.780432, 4.763298, 4.774486, 4.769708, 4.766465, 4.746224, 4.7384205, 4.733393, 4.7313013, 4.7239223, 4.7337465, 4.7348127, 4.7375097, 4.7386513, 4.7384, 4.7365046, 4.7369394, 4.738298, 4.750876, 4.749951, 4.743178, 4.738339, 4.7406154, 4.7438307, 4.7428856, 4.7427635, 4.745714, 4.7469854, 4.7456937, 4.745945, 4.747414, 4.7464075, 4.7461424, 4.7484684, 4.749067, 4.749815, 4.7514, 4.756748, 4.7530737, 4.760145, 4.766942, 4.764919, 4.7735047, 4.767371, 4.7752905, 4.7886744, 4.798904, 4.7967315, 4.781326, 4.8011794, 4.8031816, 4.7939453, 4.762399, 4.7676234, 4.787235, 4.7775064, 4.7762313, 4.774302, 4.7738247, 4.768761, 4.7673783, 4.775113, 4.7826695, 4.7721615, 4.774786, 4.7761974, 4.785317, 4.779164, 4.7809234, 4.8075633, 4.813903, 4.816154, 4.8136773, 4.827997, 4.8286753, 4.845182, 4.837659, 4.845525, 4.8435354, 4.829059, 4.817906, 4.795393, 4.7988014, 4.8020263, 4.8161607, 4.8076453, 4.80582, 4.8013844, 4.8077617, 4.8078775, 4.8366995, 4.8363566, 4.8381524, 4.827922, 4.8381734, 4.8424177, 4.855895, 4.8537736, 4.8152575, 4.8134856, 4.8156614, 4.843652, 4.81718, 4.815805, 4.816831, 4.818323, 4.8121314, 4.8116937, 4.812952, 4.815935, 4.841197, 4.8411283, 4.8422256, 4.845106, 4.844791, 4.845991, 4.8512063, 4.8259015, 4.8247237, 4.8212867, 4.848214, 4.856403, 4.819979, 4.804938, 4.804309, 4.8122473, 4.8115635, 4.8239775, 4.820089, 4.806729, 4.8024025, 4.811133, 4.8093615, 4.8097787, 4.801972, 4.782874, 4.802211, 4.8074265, 4.817112, 4.819617, 4.7859373, 4.7767286, 4.7805204, 4.7696877, 4.77527, 4.792907, 4.7930026, 4.7736545, 4.766499, 4.7589264, 4.755993, 4.740921, 4.741574, 4.743205, 4.7655864, 4.7782702, 4.7841296, 4.753713, 4.7638836, 4.76116, 4.753958, 4.752386, 4.75749, 4.775379, 4.766411, 4.7616706, 4.7592874, 4.7723117, 4.795707, 4.788374, 4.8015485, 4.786702, 4.7638087, 4.7558093, 4.75438, 4.746795, 4.7433753, 4.7494135, 4.7492027, 4.747536, 4.7495155, 4.749155, 4.73609, 4.7289996, 4.7297735, 4.7373266, 4.7423897, 4.7331624, 4.7311926, 4.7294, 4.7288094, 4.7264066, 4.7264266, 4.72568, 4.7254224, 4.7253475, 4.7262707, 4.7272615, 4.7272143, 4.726569, 4.7292237, 4.729672, 4.730351, 4.7301064, 4.730908, 4.732388, 4.7332506, 4.731349, 4.733597, 4.7348943, 4.748931, 4.7395964, 4.741078, 4.7654095, 4.762808, 4.779, 4.7627807, 4.7690544, 4.7777658, 4.7754335, 4.7689314, 4.7583413, 4.756347, 4.7543054, 4.7586884, 4.75683, 4.758423, 4.761337, 4.765096, 4.7646875, 4.7666426, 4.7779565, 4.7893705, 4.8075633, 4.8290453, 4.8264494, 4.817598, 4.824635, 4.789596, 4.7924294, 4.794908, 4.792559, 4.7807255, 4.7777996, 4.7815576, 4.78445, 4.786354, 4.79288, 4.7956934, 4.7897735, 4.788074, 4.781073, 4.7938766, 4.799068, 4.797852, 4.7827854, 4.776961, 4.787746, 4.77542, 4.7889676, 4.8105855, 4.7887907, 4.7797227, 4.772209, 4.7672215, 4.7720795, 4.768938, 4.764885, 4.7648644, 4.764973, 4.765375, 4.7568164, 4.7637267, 4.7725363, 4.7911797, 4.789814, 4.800892, 4.830593, 4.814888, 4.818193, 4.8089924, 4.787985, 4.779238, 4.773763, 4.775154, 4.7786245, 4.811119, 4.793925, 4.7843065, 4.7742267, 4.769224, 4.7419, 4.778222, 4.7711053, 4.7395687, 4.7340994, 4.7453127, 4.742267, 4.7479515, 4.747951, 4.7507606, 4.742729, 4.7449455, 4.7407584, 4.7351794, 4.7365246, 4.7450953, 4.740588, 4.7590833, 4.7469583, 4.747815, 4.7474074, 4.758239, 4.7560816, 4.7728295, 4.774479, 4.773804, 4.7749224, 4.7755084, 4.765818, 4.764919, 4.7609825, 4.7728024, 4.7769675, 4.7737293, 4.766465, 4.7547407, 4.7525635, 4.747754, 4.7516584, 4.755993, 4.753162, 4.754679, 4.753577, 4.76259, 4.762113, 4.7622495, 4.76133, 4.762808, 4.7609215, 4.763543, 4.7507334, 4.7573476, 4.760234, 4.76133, 4.763128, 4.760976, 4.763761, 4.7658796, 4.764899, 4.7625694, 4.7636523, 4.7654233, 4.7653413, 4.7654915, 4.764728, 4.8296075, 4.7675824, 4.830039, 4.788709, 4.8082266, 4.8080826, 4.7723055, 4.755122, 4.782506, 4.752659, 4.76776, 4.748298, 4.7518153, 4.7809234, 4.775918, 4.815709, 4.782752, 4.7749295, 4.781954, 4.7612348, 4.7619634, 4.753802, 4.7735863, 4.766806, 4.7717733, 4.804808, 4.820096, 4.852737, 4.772646, 4.794956, 4.764885, 4.7880807, 4.7679095, 4.7729726, 4.7686386, 4.7586474, 4.7573543, 4.7728906, 4.7803364, 4.8122134, 4.7817755, 4.7787066, 4.8035297, 4.8092656, 4.811406, 4.7944574, 4.790217, 4.786197, 4.779845, 4.7924633, 4.786033, 4.7917805, 4.78138, 4.7632365, 4.764844, 4.7860537, 4.7869477, 4.767051, 4.7661996, 4.797401, 4.774847, 4.782015, 4.7781544, 4.7671056, 4.764381, 4.763489, 4.761187, 4.7609553, 4.759873, 4.775031, 4.7758904, 4.7782903, 4.770015, 4.7668805, 4.748169, 4.760145, 4.764946, 4.7592874, 4.766854, 4.7646194, 4.741472, 4.7432804, 4.732945, 4.727146, 4.7506175, 4.728538, 4.7268405, 4.724689, 4.7130694, 4.7094088, 4.713944, 4.7196274, 4.723427, 4.719315, 4.7260127, 4.7194033, 4.727391, 4.7325444, 5.1477666, 0.03126, 0.0335193, 0.0210293, 0.0192077, 0.0182964, 0.0797143, 0.0063158, 0.0059825, 0.0057381, 0.0055825, 0.0055103, 0.0054798, 0.0054603, 0.0054882, 0.0059408, 0.0060466, 0.0060553, 0.006061, 0.0060358, 0.142353, 0.0643376, 0.0270711, 0.0537039, 0.100791, 0.1364123, 0.1502624, 0.1514896, 0.1490687, 0.1459698, 0.1429317, 0.1403186, 0.1379366, 0.1359536, 0.1343183, 0.1330239, 0.131807, 0.1308623, 0.1300744, 0.1293811, 0.1288267, 0.128181, 0.1273911, 0.1266369, 0.1259359, 0.1253765, 0.1247112, 0.1240638, 0.1233548, 0.1226784, 0.1219023, 0.1210912, 0.1203362, 0.1195756, 0.1189092, 0.1182723, 0.1176445, 0.1170461, 0.11636, 0.115677, 0.1150645, 0.1144903, 0.1139133, 0.1133423, 0.1127861, 0.1122125, 0.1115835, 0.1110015, 0.1104108, 0.1098028, 0.1091978, 0.108558, 0.1079213, 0.1073227, 0.1067068, 0.1061202, 0.1055105, 0.1049301, 0.1043353, 0.1037814, 0.103219, 0.1026305, 0.1020713, 0.1015326, 0.1009911, 0.1004905, 0.1000017, 0.0995682, 0.0991726, 0.098812, 0.098498, 0.0981928, 0.0978934, 0.097594, 0.0972744, 0.0969286, 0.0965713, 0.0961937, 0.0957959, 0.0953546, 0.0949018, 0.0944606, 0.0940341, 0.0936077, 0.0931436, 0.0927174, 0.0923144, 0.0919347, 0.0915811, 0.0912247, 0.0908973, 0.0905932, 0.0903209, 0.0900574, 0.0898171, 0.0895565, 0.0892902, 0.0890267, 0.0887489, 0.0884711, 0.0881933, 0.0879069, 0.0876119, 0.0873169, 0.0870335, 0.0867704, 0.0865218, 0.0862645, 0.0860073, 0.0857761, 0.0855507, 0.0853311, 0.0850999, 0.0848602, 0.0846031, 0.0843432, 0.084066, 0.0837715, 0.0834742, 0.0831653, 0.0828363, 0.0824959, 0.0821583, 0.0818209, 0.0814459, 0.0810567, 0.080656, 0.0802323, 0.0798, 0.0794024, 0.0012128, 0.0010795, 0.0010685, 0.0010546, 0.0010573, 0.0010712, 0.0010935, 0.0010714}
CNDC_quality_control =
  {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
PSAL =
  {35.7194, 35.7227, 35.7205, 35.7191, 35.7166, 35.7175, 35.7125, 35.7121, 35.7181, 35.7196, 35.7165, 35.717, 35.7313, 35.734, 35.7318, 35.7297, 35.7274, 35.7286, 35.7262, 35.7215, 35.7246, 35.7207, 35.7153, 35.7127, 35.7124, 35.7118, 35.7127, 35.7346, 35.7261, 35.7261, 35.724, 35.7325, 35.7374, 35.7299, 35.7287, 35.7383, 35.7419, 35.7385, 35.7348, 35.7336, 35.7403, 35.7445, 35.7425, 35.746, 35.7441, 35.7477, 35.7448, 35.748, 35.7467, 35.7465, 35.747, 35.748, 35.7473, 35.7447, 35.7474, 35.7371, 35.7366, 35.7265, 35.7326, 35.7263, 35.7275, 35.7229, 35.72, 35.7227, 35.7215, 35.7209, 35.7206, 35.7232, 35.7238, 35.7248, 35.7278, 35.7262, 35.7179, 35.7174, 35.7171, 35.7231, 35.7258, 35.7231, 35.7273, 35.7361, 35.7702, 35.7601, 35.7759, 35.775, 35.7809, 35.7846, 35.7818, 35.7844, 35.7852, 35.7869, 35.7853, 35.781, 35.7852, 35.7836, 35.7839, 35.7841, 35.7806, 35.7674, 35.7738, 35.7623, 35.7526, 35.752, 35.7528, 35.7535, 35.7541, 35.7536, 35.7534, 35.7539, 35.7495, 35.7557, 35.7555, 35.7539, 35.7526, 35.7611, 35.7497, 35.7545, 35.7542, 35.7537, 35.7558, 35.7551, 35.7552, 35.7566, 35.7564, 35.759, 35.7663, 35.76, 35.7704, 35.7745, 35.7754, 35.7821, 35.7789, 35.7794, 35.7794, 35.7736, 35.7713, 35.7703, 35.7684, 35.7658, 35.7649, 35.7634, 35.7644, 35.7613, 35.7629, 35.7675, 35.7621, 35.7619, 35.7623, 35.7587, 35.7591, 35.7605, 35.7569, 35.7599, 35.7586, 35.7541, 35.7548, 35.7562, 35.7574, 35.7526, 35.759, 35.7549, 35.7514, 35.7517, 35.7492, 35.7563, 35.7532, 35.7541, 35.7586, 35.7702, 35.7541, 35.7446, 35.7573, 35.7688, 35.7471, 35.7384, 35.7607, 35.7496, 35.7454, 35.746, 35.7738, 35.766, 35.7374, 35.7607, 35.7446, 35.7472, 35.7501, 35.7882, 35.7673, 35.7643, 35.7636, 35.7642, 35.7644, 35.7651, 35.7648, 35.7646, 35.7642, 35.7645, 35.7651, 35.765, 35.7652, 35.7654, 35.7653, 35.7648, 35.7651, 35.7645, 35.7656, 35.7651, 35.7664, 35.7628, 35.7641, 35.7639, 35.7662, 35.7667, 35.7664, 35.7598, 35.7586, 35.7707, 35.7661, 35.7637, 35.7578, 35.7582, 35.762, 35.7587, 35.7592, 35.758, 35.7525, 35.7536, 35.7531, 35.7502, 35.7539, 35.7543, 35.7615, 35.7502, 35.7583, 35.758, 35.7514, 35.7505, 35.7516, 35.7511, 35.7518, 35.7527, 35.75, 35.7543, 35.7593, 35.764, 35.7639, 35.7621, 35.7643, 35.768, 35.7688, 35.7701, 35.7646, 35.7611, 35.7664, 35.7662, 35.7662, 35.7671, 35.7654, 35.7659, 35.7635, 35.7661, 35.7647, 35.761, 35.7553, 35.764, 35.7669, 35.7638, 35.7603, 35.7598, 35.764, 35.7601, 35.7603, 35.7614, 35.7566, 35.756, 35.7646, 35.7568, 35.765, 35.7604, 35.7732, 35.7618, 35.7571, 35.7625, 35.7691, 35.7631, 35.7618, 35.7593, 35.7568, 35.7677, 35.7605, 35.7706, 35.7588, 35.7638, 35.7576, 35.761, 35.7659, 35.7579, 35.7566, 35.7576, 35.7609, 35.7583, 35.7599, 35.7585, 35.7576, 35.7536, 35.7596, 35.7601, 35.7607, 35.7554, 35.7602, 35.7606, 35.7609, 35.7575, 35.7618, 35.7608, 35.7636, 35.7606, 35.7609, 35.7585, 35.7622, 35.7625, 35.7611, 35.7588, 35.757, 35.7639, 35.7598, 35.7646, 35.7646, 35.7599, 35.7588, 35.7626, 35.7605, 35.7609, 35.7628, 35.7563, 35.7595, 35.7647, 35.7601, 35.7622, 35.7608, 35.7546, 35.7583, 35.7578, 35.758, 35.7523, 35.7597, 35.7665, 35.7605, 35.7594, 35.7668, 35.749, 35.7629, 35.7606, 35.7639, 35.7663, 35.7627, 35.764, 35.7607, 35.7664, 35.7646, 35.7658, 35.7629, 35.7617, 35.7639, 35.7687, 35.768, 35.7664, 35.767, 35.7668, 35.7698, 35.7685, 35.7691, 35.7701, 35.7631, 35.7752, 35.766, 35.7664, 35.7674, 35.7706, 35.775, 35.7727, 35.7714, 35.7748, 35.7746, 35.7739, 35.7743, 35.7707, 35.7729, 35.7708, 35.775, 35.774, 35.7705, 35.7651, 35.7686, 35.7687, 35.7675, 35.7658, 35.764, 35.769, 35.767, 35.7645, 35.7645, 35.7652, 35.766, 35.7663, 35.7644, 35.7646, 35.7648, 35.7643, 35.7651, 35.7669, 35.7654, 35.7601, 35.7665, 35.7691, 35.758, 35.7644, 35.7695, 35.7766, 35.7649, 35.7622, 35.7609, 35.7638, 35.7651, 35.7638, 35.7631, 35.7622, 35.7594, 35.7616, 35.7625, 35.7651, 35.766, 35.7594, 35.7651, 35.7592, 35.7657, 35.7656, 35.7653, 35.7628, 35.7658, 35.7603, 35.7596, 35.7629, 35.7643, 35.7619, 35.7587, 35.7599, 35.7593, 35.7621, 35.7612, 35.7611, 35.7611, 35.7594, 35.7602, 35.7606, 35.7622, 35.761, 35.7593, 35.7601, 35.7605, 35.7596, 35.7598, 35.7604, 35.7594, 35.7602, 35.7598, 35.7604, 35.7595, 35.7603, 35.759, 35.7588, 35.7583, 35.7592, 35.7603, 35.754, 35.7564, 35.7558, 35.7595, 35.754, 35.7537, 35.7599, 35.7547, 35.7536, 35.7581, 35.7584, 35.754, 35.7594, 35.7554, 35.7594, 35.7531, 35.7557, 35.7562, 35.7572, 35.7562, 35.7561, 35.7537, 35.7548, 35.7554, 35.754, 35.7547, 35.7522, 35.7545, 35.7518, 35.7428, 35.7462, 35.7476, 35.7477, 35.7361, 35.741, 35.7316, 35.7411, 35.7361, 35.7397, 35.7413, 35.7457, 35.7502, 35.7459, 35.7489, 35.7431, 35.7436, 35.7457, 35.7536, 35.7478, 35.7492, 35.7341, 35.7414, 35.7398, 35.7447, 35.7372, 35.7435, 35.7423, 35.7458, 35.7603, 35.7555, 35.7548, 35.7328, 35.7569, 35.7555, 35.755, 35.7569, 35.7616, 35.7589, 35.7584, 35.7579, 35.7474, 35.7569, 35.7518, 35.755, 35.7555, 35.7534, 35.7433, 35.7599, 35.7565, 35.7551, 35.7525, 35.7505, 35.7636, 35.759, 35.7566, 35.7571, 35.7601, 35.7615, 35.7621, 35.7581, 35.7598, 35.7578, 35.7597, 35.7604, 35.7579, 35.753, 35.7453, 35.7593, 35.7588, 35.7616, 35.7571, 35.7549, 35.7546, 35.7557, 35.7538, 35.7553, 35.7572, 35.7591, 35.7581, 35.756, 35.7522, 35.7508, 35.7523, 35.7461, 35.7537, 35.7595, 35.7546, 35.749, 35.7496, 35.7593, 35.7559, 35.7566, 35.7556, 35.7542, 35.7544, 35.7593, 35.7587, 35.7538, 35.7576, 35.7592, 35.7582, 35.7593, 35.7589, 35.7585, 35.7576, 35.7587, 35.7561, 35.7572, 35.7561, 35.7556, 35.7546, 35.7568, 35.7607, 35.7598, 35.7586, 35.7561, 35.758, 35.7596, 35.7591, 35.76, 35.7601, 35.7594, 35.7595, 35.759, 35.7596, 35.7595, 35.7594, 35.7591, 35.7596, 35.7581, 35.7585, 35.7588, 35.7592, 35.7588, 35.7592, 35.759, 35.7583, 35.7587, 35.759, 35.7589, 35.7512, 35.7635, 35.7553, 35.7556, 35.7533, 35.7534, 35.7603, 35.7567, 35.754, 35.7544, 35.7572, 35.7593, 35.7552, 35.7554, 35.7541, 35.7561, 35.7531, 35.7534, 35.7524, 35.7528, 35.7542, 35.747, 35.7507, 35.7524, 35.7507, 35.7575, 35.7495, 35.7556, 35.7604, 35.7537, 35.7575, 35.7593, 35.7607, 35.7606, 35.7596, 35.7598, 35.7606, 35.7592, 35.7593, 35.763, 35.7611, 35.7586, 35.7541, 35.762, 35.7634, 35.7615, 35.7587, 35.7577, 35.7624, 35.7537, 35.7596, 35.7646, 35.7607, 35.7598, 35.7613, 35.7572, 35.7604, 35.7608, 35.7596, 35.7607, 35.759, 35.7613, 35.7573, 35.7585, 35.7619, 35.761, 35.7629, 35.7559, 35.7633, 35.7589, 35.7639, 35.7617, 35.7607, 35.7601, 35.7586, 35.7598, 35.7574, 35.7674, 35.7596, 35.7601, 35.7617, 35.7611, 35.7568, 35.7595, 35.7622, 35.7589, 35.7579, 35.7573, 35.7601, 35.7614, 35.7617, 35.7587, 35.7591, 35.7595, 35.7593, 35.7578, 35.759, 35.7613, 35.7583, 35.7622, 35.7598, 35.7598, 35.7606, 35.7616, 35.7588, 35.7585, 35.7595, 35.7588, 35.7593, 35.7628, 35.7598, 35.7611, 35.7565, 35.7583, 35.761, 35.761, 35.7632, 35.7613, 35.7622, 35.7581, 35.7606, 35.7607, 35.7595, 35.7601, 35.7587, 35.7613, 35.7596, 35.7612, 35.7593, 35.7605, 35.7599, 35.7615, 35.7581, 35.7587, 35.7608, 35.7588, 35.7613, 35.7596, 35.7606, 35.7601, 35.7607, 35.7598, 35.7605, 35.759, 35.7616, 35.7574, 35.7589, 35.7626, 35.7551, 35.7804, 35.7606, 35.7361, 35.7854, 35.7614, 35.7513, 35.765, 35.7582, 35.7625, 35.7585, 35.7541, 35.7749, 35.7399, 35.7881, 35.7568, 35.7732, 35.7606, 35.7567, 35.7623, 35.7524, 35.7613, 35.7538, 35.7475, 35.742, 35.7351, 35.7685, 35.7582, 35.7652, 35.7454, 35.7537, 35.7467, 35.7537, 35.7538, 35.7514, 35.7381, 35.748, 35.7382, 35.7423, 35.7457, 35.7391, 35.7528, 35.7434, 35.7537, 35.7467, 35.7572, 35.7502, 35.7579, 35.757, 35.7606, 35.7619, 35.7523, 35.7562, 35.754, 35.7598, 35.7626, 35.7623, 35.7581, 35.7598, 35.7725, 35.7682, 35.761, 35.7609, 35.7625, 35.7607, 35.7603, 35.7581, 35.7568, 35.7577, 35.753, 35.7633, 35.7611, 35.767, 35.7645, 35.7637, 35.7639, 35.7627, 35.7592, 35.7618, 35.77, 35.7553, 35.7543, 35.7544, 35.7523, 35.7478, 35.7442, 35.746, 35.7458, 35.7448, 35.7464, 35.7481, 35.7528, 35.7523, 35.7558, 35.757, 35.757, 35.6399, 0.1511, 0.1702, 0.1041, 0.0975, 0.093, 0.3949, 0.0364, 0.0349, 0.0339, 0.0332, 0.0329, 0.0327, 0.0326, 0.0327, 0.0348, 0.0351, 0.0349, 0.0347, 0.0348, 0.6783, 0.2949, 0.1241, 0.2458, 0.4693, 0.6432, 0.7122, 0.7189, 0.7076, 0.693, 0.6787, 0.6666, 0.6557, 0.6468, 0.6397, 0.6342, 0.6291, 0.6253, 0.6224, 0.6198, 0.618, 0.6157, 0.6126, 0.6097, 0.6071, 0.6052, 0.6027, 0.6003, 0.5976, 0.5952, 0.5921, 0.5888, 0.5859, 0.5831, 0.5807, 0.5783, 0.5762, 0.5741, 0.5714, 0.5689, 0.5666, 0.5645, 0.5624, 0.5603, 0.5582, 0.5561, 0.5536, 0.5514, 0.549, 0.5465, 0.5441, 0.5415, 0.5388, 0.5364, 0.5338, 0.5314, 0.5289, 0.5267, 0.5243, 0.5222, 0.5201, 0.5179, 0.5158, 0.5137, 0.5116, 0.5096, 0.5076, 0.5059, 0.5042, 0.5028, 0.5017, 0.5006, 0.4995, 0.4986, 0.4974, 0.4962, 0.4949, 0.4936, 0.492, 0.4902, 0.4885, 0.4867, 0.4851, 0.4834, 0.4815, 0.4799, 0.4782, 0.4768, 0.4755, 0.4741, 0.4729, 0.4719, 0.471, 0.4702, 0.4695, 0.4686, 0.4677, 0.4668, 0.4658, 0.4648, 0.4638, 0.4627, 0.4615, 0.4603, 0.4592, 0.4581, 0.4572, 0.4561, 0.455, 0.454, 0.4531, 0.4522, 0.4511, 0.45, 0.4487, 0.4474, 0.446, 0.4444, 0.4428, 0.4411, 0.4393, 0.4373, 0.4354, 0.4334, 0.4312, 0.429, 0.4266, 0.4241, 0.4216, 0.4192, 0.0147, 0.014, 0.014, 0.0139, 0.0139, 0.014, 0.0141, 0.0141}
PSAL_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {81.291, 81.001, 81.037, 81.069, 81.171, 81.1, 81.082, 81.093, 81.0, 81.045, 81.243, 81.044, 81.012, 81.202, 80.958, 81.185, 81.11, 80.965, 81.187, 81.148, 80.977, 81.257, 81.187, 81.238, 81.269, 81.295, 81.202, 81.041, 81.177, 81.106, 81.14, 81.066, 81.167, 81.225, 81.289, 81.263, 81.333, 81.342, 81.275, 81.268, 81.255, 81.404, 81.335, 81.169, 81.38, 81.245, 81.287, 81.238, 81.315, 81.179, 81.368, 81.355, 81.39, 81.446, 81.287, 81.367, 81.239, 81.159, 81.341, 81.315, 81.226, 81.25, 81.416, 81.335, 81.28, 81.428, 81.26, 81.288, 81.309, 81.286, 81.362, 81.322, 81.368, 81.429, 81.359, 81.432, 81.414, 81.172, 81.389, 81.312, 81.234, 81.207, 81.38, 81.346, 81.172, 81.365, 81.173, 81.282, 81.219, 81.272, 81.201, 81.28, 81.313, 81.288, 81.331, 81.208, 81.105, 81.155, 81.096, 81.051, 81.06, 81.072, 81.176, 81.0, 80.938, 81.236, 81.044, 81.154, 81.043, 81.073, 81.127, 81.204, 81.245, 81.103, 81.086, 81.059, 81.073, 80.962, 80.966, 81.025, 80.997, 81.029, 80.975, 81.031, 80.891, 80.993, 80.896, 81.031, 81.07, 80.847, 81.072, 80.884, 81.081, 80.989, 80.824, 80.82, 80.859, 80.764, 80.962, 80.922, 80.792, 80.96, 80.857, 80.92, 80.948, 80.965, 80.835, 80.954, 80.878, 81.024, 81.104, 80.999, 80.984, 80.95, 81.007, 80.883, 80.977, 80.988, 81.011, 80.99, 81.062, 81.059, 81.151, 81.014, 81.084, 80.929, 81.056, 81.091, 81.204, 81.003, 81.053, 81.092, 81.11, 81.148, 81.012, 81.171, 81.094, 80.997, 80.983, 81.093, 81.298, 81.166, 81.135, 81.289, 81.153, 81.096, 81.206, 81.27, 81.14, 81.159, 81.058, 81.254, 81.316, 81.175, 81.192, 81.283, 81.236, 81.219, 81.338, 81.28, 81.36, 81.232, 81.198, 81.389, 81.355, 81.322, 81.251, 81.231, 81.337, 81.374, 81.336, 81.226, 81.355, 81.395, 81.252, 81.327, 81.227, 81.415, 81.224, 81.301, 81.307, 81.271, 81.142, 81.178, 81.201, 81.227, 81.151, 81.27, 81.276, 81.164, 81.194, 81.097, 81.383, 81.037, 81.251, 81.203, 81.105, 81.147, 81.128, 81.106, 81.032, 81.021, 80.938, 81.085, 81.045, 80.915, 80.924, 80.948, 81.006, 80.924, 81.196, 80.981, 80.847, 80.883, 81.114, 80.978, 80.731, 80.854, 81.049, 80.884, 81.011, 80.899, 80.986, 80.781, 80.865, 80.798, 80.831, 80.913, 80.856, 80.884, 80.832, 80.996, 80.933, 80.934, 80.874, 80.986, 80.837, 81.058, 80.805, 80.68, 80.913, 80.891, 80.935, 80.79, 80.878, 80.866, 80.841, 80.905, 80.907, 81.06, 80.849, 80.88, 80.911, 80.986, 80.897, 80.913, 81.001, 80.903, 80.942, 81.093, 80.963, 80.867, 80.988, 81.117, 81.122, 81.015, 81.018, 81.17, 81.074, 81.03, 81.031, 81.175, 80.978, 80.762, 81.027, 81.126, 81.141, 81.033, 81.147, 81.068, 81.045, 81.301, 81.259, 80.995, 81.185, 81.197, 81.061, 81.246, 81.208, 81.076, 81.262, 81.252, 81.191, 81.328, 81.283, 81.191, 81.287, 81.233, 81.343, 81.325, 81.452, 81.343, 81.463, 81.376, 81.371, 81.287, 81.452, 81.457, 81.471, 81.487, 81.356, 81.487, 81.417, 81.516, 81.262, 81.415, 81.438, 81.413, 81.31, 81.31, 81.335, 81.488, 81.416, 81.52, 81.544, 81.2, 81.257, 81.281, 81.523, 81.288, 81.244, 81.324, 81.347, 81.256, 81.329, 81.289, 81.518, 81.383, 81.155, 81.261, 81.242, 81.184, 81.131, 81.208, 81.055, 81.206, 81.133, 81.215, 81.051, 81.114, 81.075, 81.117, 80.874, 81.145, 81.033, 80.95, 80.975, 81.003, 81.092, 80.97, 80.904, 81.017, 80.749, 80.92, 80.917, 80.753, 80.64, 80.98, 80.92, 80.812, 80.688, 80.989, 80.709, 80.728, 80.942, 81.051, 80.959, 80.868, 80.722, 80.944, 80.914, 80.796, 80.755, 80.909, 80.775, 80.825, 80.956, 80.813, 80.93, 80.85, 80.849, 80.677, 80.787, 80.938, 80.849, 80.875, 80.938, 80.878, 80.837, 80.824, 80.852, 81.072, 81.029, 80.913, 81.048, 81.044, 80.935, 81.02, 81.026, 81.019, 81.118, 81.003, 81.129, 81.073, 81.001, 81.154, 81.09, 81.064, 81.127, 81.271, 81.07, 81.193, 81.103, 81.274, 80.963, 81.262, 81.039, 81.22, 81.13, 81.165, 81.09, 81.062, 81.209, 81.218, 81.397, 81.329, 81.202, 81.22, 81.273, 81.155, 81.271, 81.183, 81.411, 81.462, 81.321, 81.35, 81.456, 81.595, 81.495, 81.297, 81.303, 81.443, 81.578, 81.537, 81.51, 81.325, 81.373, 81.55, 81.5, 81.725, 81.484, 81.494, 81.726, 81.488, 81.428, 81.615, 81.646, 81.443, 81.517, 81.371, 81.537, 81.526, 81.471, 81.434, 81.549, 81.449, 81.34, 81.359, 81.549, 81.334, 81.52, 81.56, 81.337, 81.452, 81.354, 81.187, 81.283, 81.426, 81.109, 81.201, 81.2, 81.081, 81.196, 81.124, 81.165, 81.087, 81.135, 81.088, 80.996, 81.152, 81.042, 81.063, 80.88, 80.924, 80.763, 81.06, 80.757, 80.854, 80.786, 80.902, 80.782, 80.6, 80.832, 81.099, 80.867, 80.691, 80.933, 80.792, 80.899, 80.817, 80.787, 80.904, 80.662, 80.807, 81.006, 80.685, 80.861, 80.924, 80.715, 80.916, 80.947, 80.901, 80.942, 80.671, 80.682, 80.771, 80.887, 80.945, 80.841, 80.915, 80.999, 81.03, 80.97, 80.954, 80.965, 80.896, 80.986, 81.115, 81.133, 81.233, 81.254, 81.172, 81.218, 81.072, 81.002, 81.164, 81.228, 81.014, 81.177, 81.329, 81.102, 81.201, 81.033, 81.218, 81.062, 81.127, 80.951, 81.135, 81.201, 81.227, 81.081, 81.134, 81.149, 81.104, 81.276, 81.395, 81.493, 81.263, 81.394, 81.293, 81.344, 81.31, 81.391, 81.181, 81.307, 81.121, 81.356, 81.248, 81.563, 81.307, 81.333, 81.371, 81.318, 81.406, 81.27, 81.279, 81.304, 81.421, 81.431, 81.311, 81.494, 81.384, 81.536, 81.307, 81.478, 81.449, 81.518, 81.468, 81.63, 81.522, 81.532, 81.447, 81.425, 81.481, 81.553, 81.557, 81.331, 81.443, 81.467, 81.385, 81.428, 81.508, 81.419, 81.598, 81.489, 81.392, 81.482, 81.475, 81.459, 81.421, 81.251, 81.24, 81.384, 81.114, 81.204, 81.213, 81.298, 81.289, 81.054, 81.024, 81.169, 81.143, 81.024, 81.392, 81.032, 81.041, 80.914, 80.893, 81.012, 80.856, 80.775, 80.95, 80.948, 80.921, 80.924, 80.873, 80.817, 80.796, 80.806, 80.957, 80.805, 80.739, 80.716, 80.743, 80.755, 80.812, 80.84, 80.816, 80.672, 80.77, 80.656, 80.722, 80.984, 80.706, 80.728, 80.623, 80.63, 80.641, 80.953, 80.978, 80.885, 80.774, 80.744, 80.986, 80.836, 81.08, 80.868, 80.84, 80.995, 80.982, 80.769, 80.981, 80.812, 81.026, 80.978, 81.015, 81.026, 81.118, 81.098, 81.062, 80.903, 81.118, 81.001, 81.057, 81.094, 81.001, 81.069, 81.088, 80.991, 81.153, 81.062, 81.073, 81.027, 80.935, 81.019, 81.081, 81.148, 81.108, 81.025, 81.038, 81.13, 81.118, 81.099, 81.209, 81.184, 81.07, 81.16, 81.224, 81.248, 81.182, 81.137, 81.177, 81.286, 81.195, 81.237, 81.256, 81.219, 81.303, 81.341, 81.25, 81.293, 81.309, 81.321, 81.395, 81.338, 81.344, 81.401, 81.484, 81.438, 81.644, 81.342, 81.651, 81.475, 81.62, 81.429, 81.499, 81.48, 81.56, 81.433, 81.522, 81.537, 81.595, 81.65, 81.572, 81.586, 81.605, 81.512, 81.691, 81.428, 81.597, 81.572, 81.629, 81.547, 81.5, 81.63, 81.675, 81.59, 81.24, 81.559, 81.317, 81.477, 81.289, 81.395, 81.3, 81.194, 81.338, 81.249, 81.202, 81.294, 81.116, 81.161, 81.279, 81.1, 81.146, 81.216, 81.054, 81.13, 80.997, 81.029, 80.926, 81.029, 80.774, 80.857, 81.027, 81.012, 80.975, 80.954, 80.819, 80.897, 80.823, 80.889, 80.881, 80.819, 80.849, 80.933, 80.924, 80.793, 80.917, 80.909, 81.09, 80.908, 81.031, 80.994, 80.865, 80.951, 81.07, 81.096, 81.208, 81.023, 80.954, 81.267, 81.023, 81.019, 81.293, 81.124, 81.194, 81.171, 81.282, 81.318, 81.435, 81.35, 81.489, 81.285, 81.62, 81.294, 81.411, 81.464, 3.165, 1.94, 0.007, -0.027, -0.028, -0.025, 0.069, -0.016, -0.017, -0.017, -0.021, -0.02, -0.021, -0.022, -0.026, -0.028, -0.028, -0.035, -0.041, -0.058, 0.109, 0.091, 0.085, 0.128, 0.134, 0.134, 0.134, 0.132, 0.131, 0.129, 0.13, 0.129, 0.129, 0.129, 0.126, 0.125, 0.126, 0.124, 0.123, 0.124, 0.123, 0.124, 0.124, 0.125, 0.126, 0.126, 0.128, 0.129, 0.127, 0.128, 0.13, 0.128, 0.129, 0.13, 0.131, 0.133, 0.135, 0.133, 0.136, 0.135, 0.134, 0.134, 0.135, 0.136, 0.137, 0.137, 0.137, 0.134, 0.137, 0.136, 0.139, 0.136, 0.134, 0.135, 0.136, 0.136, 0.136, 0.138, 0.137, 0.138, 0.138, 0.139, 0.141, 0.14, 0.14, 0.142, 0.14, 0.14, 0.139, 0.138, 0.14, 0.14, 0.136, 0.139, 0.138, 0.138, 0.137, 0.137, 0.138, 0.137, 0.138, 0.137, 0.138, 0.139, 0.138, 0.142, 0.142, 0.142, 0.143, 0.146, 0.146, 0.147, 0.145, 0.147, 0.147, 0.145, 0.147, 0.146, 0.148, 0.149, 0.149, 0.149, 0.15, 0.15, 0.152, 0.155, 0.154, 0.158, 0.157, 0.156, 0.157, 0.156, 0.156, 0.155, 0.157, 0.157, 0.155, 0.155, 0.155, 0.159, 0.16, 0.161, 0.16, 0.16, 0.159, 0.159, 0.16, 0.162, 0.159, 0.162, 0.005, -0.038, -0.036, -0.046, -0.069, -0.033, -0.033, -0.033}
PRES_REL_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {80.708, 80.421, 80.457, 80.489, 80.59, 80.52, 80.502, 80.512, 80.42, 80.465, 80.661, 80.464, 80.432, 80.62, 80.378, 80.604, 80.529, 80.385, 80.605, 80.567, 80.397, 80.675, 80.605, 80.656, 80.687, 80.713, 80.62, 80.46, 80.596, 80.525, 80.559, 80.485, 80.586, 80.643, 80.707, 80.681, 80.75, 80.759, 80.693, 80.686, 80.673, 80.821, 80.752, 80.587, 80.797, 80.663, 80.705, 80.656, 80.732, 80.598, 80.786, 80.772, 80.807, 80.863, 80.705, 80.784, 80.657, 80.578, 80.758, 80.732, 80.644, 80.668, 80.833, 80.752, 80.698, 80.845, 80.677, 80.706, 80.726, 80.704, 80.78, 80.739, 80.786, 80.846, 80.776, 80.849, 80.831, 80.591, 80.806, 80.73, 80.653, 80.625, 80.797, 80.763, 80.591, 80.782, 80.592, 80.7, 80.637, 80.689, 80.619, 80.698, 80.731, 80.706, 80.749, 80.626, 80.524, 80.574, 80.515, 80.471, 80.479, 80.491, 80.594, 80.42, 80.358, 80.654, 80.464, 80.573, 80.462, 80.492, 80.546, 80.623, 80.663, 80.522, 80.505, 80.478, 80.492, 80.382, 80.386, 80.445, 80.417, 80.448, 80.395, 80.451, 80.312, 80.413, 80.316, 80.451, 80.49, 80.268, 80.491, 80.305, 80.5, 80.409, 80.245, 80.242, 80.28, 80.186, 80.382, 80.343, 80.213, 80.381, 80.278, 80.34, 80.369, 80.385, 80.256, 80.375, 80.299, 80.443, 80.523, 80.419, 80.404, 80.37, 80.427, 80.303, 80.397, 80.408, 80.43, 80.41, 80.481, 80.478, 80.569, 80.434, 80.503, 80.35, 80.476, 80.51, 80.623, 80.423, 80.472, 80.511, 80.529, 80.567, 80.432, 80.59, 80.514, 80.417, 80.403, 80.512, 80.715, 80.585, 80.554, 80.707, 80.572, 80.515, 80.624, 80.688, 80.559, 80.578, 80.478, 80.672, 80.733, 80.593, 80.611, 80.701, 80.654, 80.637, 80.756, 80.698, 80.777, 80.65, 80.617, 80.806, 80.772, 80.739, 80.669, 80.649, 80.755, 80.791, 80.753, 80.644, 80.772, 80.812, 80.67, 80.744, 80.645, 80.832, 80.642, 80.719, 80.725, 80.689, 80.561, 80.597, 80.619, 80.645, 80.569, 80.688, 80.694, 80.582, 80.612, 80.516, 80.8, 80.457, 80.669, 80.622, 80.524, 80.566, 80.547, 80.525, 80.452, 80.441, 80.358, 80.504, 80.465, 80.335, 80.345, 80.369, 80.426, 80.345, 80.614, 80.401, 80.268, 80.303, 80.533, 80.398, 80.152, 80.275, 80.468, 80.305, 80.43, 80.32, 80.405, 80.202, 80.286, 80.219, 80.252, 80.333, 80.277, 80.305, 80.253, 80.416, 80.353, 80.354, 80.295, 80.405, 80.258, 80.478, 80.226, 80.103, 80.333, 80.312, 80.356, 80.212, 80.299, 80.287, 80.262, 80.326, 80.327, 80.479, 80.27, 80.301, 80.332, 80.405, 80.318, 80.333, 80.421, 80.324, 80.363, 80.512, 80.383, 80.288, 80.408, 80.536, 80.541, 80.435, 80.438, 80.588, 80.493, 80.449, 80.451, 80.593, 80.398, 80.183, 80.447, 80.544, 80.56, 80.453, 80.566, 80.487, 80.465, 80.719, 80.677, 80.415, 80.604, 80.616, 80.48, 80.664, 80.626, 80.496, 80.68, 80.67, 80.61, 80.745, 80.701, 80.61, 80.705, 80.651, 80.761, 80.743, 80.869, 80.761, 80.879, 80.793, 80.788, 80.705, 80.869, 80.873, 80.888, 80.903, 80.774, 80.903, 80.834, 80.932, 80.68, 80.832, 80.854, 80.829, 80.727, 80.727, 80.752, 80.904, 80.833, 80.936, 80.96, 80.618, 80.675, 80.699, 80.939, 80.706, 80.662, 80.742, 80.764, 80.674, 80.746, 80.707, 80.934, 80.8, 80.574, 80.679, 80.66, 80.603, 80.55, 80.626, 80.474, 80.624, 80.552, 80.634, 80.471, 80.533, 80.495, 80.536, 80.295, 80.563, 80.453, 80.37, 80.395, 80.423, 80.511, 80.39, 80.325, 80.436, 80.17, 80.34, 80.338, 80.175, 80.062, 80.4, 80.34, 80.233, 80.11, 80.409, 80.131, 80.15, 80.363, 80.471, 80.379, 80.289, 80.144, 80.364, 80.334, 80.218, 80.176, 80.329, 80.196, 80.246, 80.376, 80.234, 80.351, 80.271, 80.27, 80.099, 80.208, 80.358, 80.27, 80.296, 80.358, 80.299, 80.258, 80.245, 80.272, 80.491, 80.448, 80.333, 80.467, 80.464, 80.356, 80.44, 80.446, 80.439, 80.537, 80.423, 80.548, 80.492, 80.421, 80.573, 80.509, 80.484, 80.546, 80.689, 80.49, 80.611, 80.522, 80.692, 80.383, 80.68, 80.459, 80.638, 80.549, 80.584, 80.509, 80.481, 80.628, 80.636, 80.814, 80.746, 80.62, 80.638, 80.691, 80.574, 80.689, 80.601, 80.828, 80.878, 80.738, 80.768, 80.872, 81.01, 80.911, 80.714, 80.72, 80.859, 80.993, 80.953, 80.926, 80.743, 80.79, 80.966, 80.916, 81.139, 80.901, 80.91, 81.141, 80.904, 80.845, 81.03, 81.061, 80.859, 80.933, 80.788, 80.953, 80.942, 80.888, 80.851, 80.965, 80.865, 80.757, 80.776, 80.965, 80.751, 80.936, 80.976, 80.755, 80.869, 80.771, 80.605, 80.701, 80.843, 80.528, 80.619, 80.618, 80.5, 80.614, 80.543, 80.584, 80.506, 80.554, 80.508, 80.416, 80.571, 80.461, 80.483, 80.301, 80.345, 80.185, 80.479, 80.179, 80.275, 80.207, 80.322, 80.204, 80.023, 80.253, 80.518, 80.288, 80.113, 80.353, 80.213, 80.32, 80.238, 80.208, 80.325, 80.085, 80.228, 80.426, 80.107, 80.282, 80.345, 80.137, 80.337, 80.367, 80.321, 80.363, 80.093, 80.104, 80.193, 80.308, 80.365, 80.262, 80.335, 80.419, 80.449, 80.39, 80.375, 80.385, 80.316, 80.405, 80.534, 80.552, 80.651, 80.672, 80.591, 80.636, 80.491, 80.422, 80.582, 80.647, 80.434, 80.595, 80.746, 80.521, 80.619, 80.453, 80.636, 80.481, 80.546, 80.371, 80.554, 80.619, 80.645, 80.5, 80.553, 80.568, 80.523, 80.694, 80.812, 80.909, 80.681, 80.81, 80.711, 80.762, 80.727, 80.808, 80.599, 80.725, 80.54, 80.774, 80.666, 80.979, 80.725, 80.75, 80.788, 80.736, 80.822, 80.688, 80.696, 80.721, 80.838, 80.847, 80.729, 80.91, 80.801, 80.952, 80.725, 80.895, 80.865, 80.934, 80.884, 81.046, 80.938, 80.948, 80.864, 80.841, 80.897, 80.968, 80.973, 80.749, 80.859, 80.883, 80.802, 80.845, 80.924, 80.835, 81.014, 80.905, 80.809, 80.898, 80.891, 80.876, 80.838, 80.669, 80.658, 80.801, 80.533, 80.623, 80.631, 80.715, 80.707, 80.473, 80.443, 80.587, 80.562, 80.443, 80.809, 80.452, 80.46, 80.334, 80.314, 80.432, 80.277, 80.196, 80.37, 80.369, 80.341, 80.345, 80.294, 80.238, 80.218, 80.227, 80.377, 80.226, 80.161, 80.138, 80.164, 80.176, 80.233, 80.261, 80.237, 80.094, 80.192, 80.079, 80.144, 80.404, 80.128, 80.15, 80.046, 80.053, 80.063, 80.373, 80.398, 80.306, 80.195, 80.166, 80.405, 80.257, 80.499, 80.289, 80.261, 80.415, 80.402, 80.191, 80.401, 80.233, 80.446, 80.398, 80.435, 80.446, 80.537, 80.517, 80.481, 80.324, 80.537, 80.421, 80.477, 80.514, 80.421, 80.489, 80.508, 80.411, 80.572, 80.481, 80.492, 80.447, 80.356, 80.439, 80.5, 80.567, 80.527, 80.445, 80.458, 80.549, 80.537, 80.518, 80.628, 80.603, 80.49, 80.579, 80.642, 80.666, 80.6, 80.556, 80.595, 80.704, 80.613, 80.655, 80.674, 80.637, 80.72, 80.758, 80.668, 80.711, 80.726, 80.738, 80.812, 80.756, 80.762, 80.818, 80.901, 80.854, 81.059, 80.759, 81.066, 80.891, 81.035, 80.846, 80.915, 80.896, 80.976, 80.85, 80.938, 80.953, 81.01, 81.065, 80.987, 81.002, 81.021, 80.928, 81.106, 80.845, 81.012, 80.987, 81.044, 80.962, 80.916, 81.046, 81.09, 81.005, 80.658, 80.974, 80.734, 80.894, 80.707, 80.812, 80.718, 80.612, 80.756, 80.667, 80.62, 80.712, 80.535, 80.58, 80.696, 80.519, 80.565, 80.635, 80.473, 80.549, 80.417, 80.448, 80.346, 80.448, 80.195, 80.278, 80.447, 80.432, 80.395, 80.375, 80.24, 80.318, 80.244, 80.309, 80.302, 80.24, 80.27, 80.353, 80.345, 80.214, 80.338, 80.329, 80.509, 80.328, 80.451, 80.414, 80.286, 80.371, 80.49, 80.515, 80.626, 80.442, 80.375, 80.685, 80.442, 80.439, 80.711, 80.543, 80.612, 80.59, 80.7, 80.736, 80.852, 80.768, 80.906, 80.702, 81.035, 80.712, 80.828, 80.881, 3.143, 1.927, 0.007, -0.027, -0.028, -0.025, 0.068, -0.016, -0.017, -0.017, -0.021, -0.02, -0.021, -0.022, -0.026, -0.028, -0.028, -0.034, -0.041, -0.057, 0.108, 0.09, 0.084, 0.127, 0.133, 0.133, 0.133, 0.131, 0.131, 0.128, 0.129, 0.128, 0.128, 0.128, 0.125, 0.124, 0.125, 0.124, 0.122, 0.123, 0.122, 0.123, 0.123, 0.124, 0.125, 0.125, 0.127, 0.128, 0.126, 0.127, 0.129, 0.127, 0.128, 0.129, 0.13, 0.132, 0.134, 0.132, 0.135, 0.134, 0.133, 0.133, 0.134, 0.135, 0.136, 0.136, 0.136, 0.133, 0.136, 0.135, 0.138, 0.135, 0.133, 0.134, 0.135, 0.135, 0.135, 0.137, 0.136, 0.137, 0.137, 0.138, 0.14, 0.139, 0.139, 0.141, 0.139, 0.139, 0.138, 0.137, 0.139, 0.139, 0.135, 0.138, 0.137, 0.137, 0.136, 0.136, 0.137, 0.136, 0.137, 0.136, 0.137, 0.138, 0.137, 0.141, 0.141, 0.141, 0.142, 0.145, 0.145, 0.146, 0.144, 0.146, 0.146, 0.144, 0.145, 0.145, 0.147, 0.148, 0.148, 0.148, 0.149, 0.149, 0.151, 0.153, 0.153, 0.157, 0.156, 0.154, 0.156, 0.154, 0.154, 0.154, 0.156, 0.156, 0.154, 0.154, 0.154, 0.158, 0.159, 0.16, 0.159, 0.159, 0.158, 0.158, 0.159, 0.16, 0.158, 0.16, 0.005, -0.038, -0.035, -0.045, -0.068, -0.033, -0.033, -0.033}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
