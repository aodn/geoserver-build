netcdf file-124.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (18 currently)
  variables:
    float LATITUDE(DEPTH=18);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=18);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=18);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=18);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=18);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=18);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185, 22988.187997685185}
TEMP =
  {32.1551, 32.1416, 32.1051, 32.0301, 31.9972, 31.9816, 31.9649, 31.9547, 31.9525, 31.9481, 31.9427, 31.9407, 31.9379, 31.9348, 31.9311, 31.9288, 31.9279, 31.9278}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879, 21.873, 22.867}
}
