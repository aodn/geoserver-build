netcdf file-85.nc {
  dimensions:
    DEPTH = 21;
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926, 23178.503113425926}
TEMP =
  {27.0666, 27.1102, 27.1045, 27.1025, 27.1036, 27.1039, 27.1043, 27.1052, 27.105, 27.1025, 27.0935, 27.0844, 27.0748, 27.0647, 27.0557, 27.0454, 27.0414, 27.0406, 27.0399, 27.0398, 27.0382}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.963, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872}
}
