netcdf file-105.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887, 22659.147013888887}
TEMP =
  {31.5442, 31.546, 31.5437, 31.5439, 31.5456, 31.5457, 31.5466, 31.547, 31.546, 31.5452, 31.5419, 31.5334, 31.5259, 31.5205, 31.5137, 31.5113, 31.509, 31.5065, 31.504, 31.5024, 31.5012}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89, 19.885, 20.879}
}
