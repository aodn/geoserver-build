netcdf file-4.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (48 currently)
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518, 21809.350393518518}
TEMP =
  {15.9466, 15.9615, 15.9553, 15.9497, 15.9434, 15.9374, 15.9329, 15.9294, 15.925, 15.9213, 15.9188, 15.9169, 15.9156, 15.9142, 15.9125, 15.91, 15.907, 15.9053, 15.9033, 15.9002, 15.8983, 15.8972, 15.8966, 15.897, 15.8968, 15.8958, 15.8956, 15.8952, 15.8954, 15.8963, 15.8973, 15.8956, 15.894, 15.8922, 15.8927, 15.8912, 15.8897, 15.8891, 15.8889, 15.8886, 15.8882, 15.8881, 15.888, 15.8875, 15.8863, 15.8845, 15.8847, 15.8836}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
