netcdf file-111.nc {
  dimensions:
    DEPTH = 22;
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185, 22987.73091435185}
TEMP =
  {31.9476, 31.9477, 31.944, 31.9407, 31.9399, 31.9401, 31.9404, 31.9423, 31.944, 31.9465, 31.9486, 31.949, 31.9465, 31.9455, 31.9457, 31.9434, 31.9414, 31.9399, 31.939, 31.9379, 31.9362, 31.9351}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.943, 10.936, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879, 21.872, 22.867}
}
