netcdf file-99.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (22 currently)
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668, 22658.896979166668}
TEMP =
  {31.4331, 31.4326, 31.4368, 31.4379, 31.442, 31.4453, 31.4454, 31.4458, 31.4462, 31.4462, 31.4454, 31.4461, 31.4489, 31.4511, 31.4526, 31.4538, 31.4548, 31.4559, 31.4566, 31.4572, 31.4583, 31.4603}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.995, 1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89, 19.885, 20.879, 21.873}
}
