netcdf file-53.nc {
  dimensions:
    DEPTH = 45;
  variables:
    float LATITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=45);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=45);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084}
LONGITUDE =
  {115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334}
TIME =
  {22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483, 22975.146481481483}
TEMP =
  {20.4148, 20.3521, 20.174, 20.0566, 20.0221, 20.0038, 19.9891, 19.9729, 19.9612, 19.9561, 19.9483, 19.9388, 19.9296, 19.9057, 19.8434, 19.7832, 19.7456, 19.7079, 19.6489, 19.6214, 19.5876, 19.5424, 19.5119, 19.4795, 19.4212, 19.3827, 19.3735, 19.3539, 19.3247, 19.26, 19.2089, 19.1795, 19.1367, 19.1084, 19.0884, 19.0808, 19.0795, 19.0752, 19.0756, 19.0713, 19.0715, 19.0702, 19.0716, 19.0721, 19.0698}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
