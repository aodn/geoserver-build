netcdf file-36.nc {
  dimensions:
    DEPTH = 48;
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223, 22263.120659722223}
TEMP =
  {20.8891, 20.8816, 20.8835, 20.8865, 20.883, 20.8771, 20.8692, 20.8673, 20.8664, 20.8683, 20.8695, 20.8702, 20.8742, 20.8716, 20.8576, 20.8515, 20.8466, 20.8445, 20.8436, 20.8456, 20.8432, 20.8381, 20.8319, 20.8342, 20.8399, 20.8354, 20.8335, 20.832, 20.8303, 20.8304, 20.831, 20.8318, 20.8328, 20.833, 20.8326, 20.8319, 20.8318, 20.8321, 20.8328, 20.8329, 20.8332, 20.8344, 20.8349, 20.8354, 20.8361, 20.8365, 20.8369, 20.8378}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
