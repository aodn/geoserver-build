netcdf file-1.nc {
  dimensions:
    DEPTH = 46;
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963, 21604.38619212963}
TEMP =
  {20.6617, 20.6652, 20.6659, 20.6667, 20.6672, 20.6675, 20.6676, 20.6678, 20.6683, 20.6688, 20.6693, 20.67, 20.6705, 20.671, 20.6711, 20.6712, 20.6712, 20.6713, 20.6716, 20.6719, 20.6721, 20.6721, 20.6717, 20.6707, 20.6697, 20.6693, 20.6691, 20.669, 20.6692, 20.6693, 20.6695, 20.6698, 20.6701, 20.6703, 20.6704, 20.6706, 20.6708, 20.6711, 20.6713, 20.6715, 20.6716, 20.6719, 20.6721, 20.6722, 20.6724, 20.6726}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
