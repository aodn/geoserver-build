netcdf file-130.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (27 currently)
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391}
TIME =
  {23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594, 23116.072280092594}
TEMP =
  {26.3667, 26.3718, 26.3654, 26.355, 26.3464, 26.3393, 26.3318, 26.328, 26.3269, 26.3243, 26.3188, 26.3152, 26.3128, 26.3091, 26.3084, 26.3087, 26.3089, 26.3087, 26.308, 26.3059, 26.3032, 26.302, 26.3018, 26.3012, 26.3003, 26.2999, 26.2999}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835}
}
