netcdf file-109.nc {
  dimensions:
    DEPTH = 19;
  variables:
    float LATITUDE(DEPTH=19);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=19);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=19);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=19);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=19);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=19);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926, 22752.03707175926}
TEMP =
  {30.0493, 30.052, 30.0501, 30.0527, 30.0887, 30.1304, 30.1227, 30.1097, 30.0964, 30.0875, 30.0831, 30.0798, 30.0776, 30.0766, 30.0757, 30.0748, 30.0747, 30.0747, 30.0746}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.89}
}
