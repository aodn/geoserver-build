netcdf file-56.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (47 currently)
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001, -32.001}
LONGITUDE =
  {115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166, 115.4166}
TIME =
  {23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741, 23062.22365740741}
TEMP =
  {23.2199, 23.1165, 22.9933, 22.9719, 22.9618, 22.9318, 22.9136, 22.9066, 22.9168, 22.9166, 22.9209, 22.9065, 22.8974, 22.8878, 22.8669, 22.8177, 22.7488, 22.709, 22.6676, 22.546, 22.436, 22.3638, 22.3151, 22.276, 22.267, 22.2614, 22.2628, 22.2608, 22.2608, 22.2621, 22.2612, 22.2619, 22.2617, 22.2632, 22.2627, 22.2627, 22.2631, 22.2628, 22.2636, 22.263, 22.2632, 22.2638, 22.2632, 22.2632, 22.2632, 22.2643, 22.2669}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
