netcdf file-22.nc {
  dimensions:
    DEPTH = 42;
  variables:
    float LATITUDE(DEPTH=42);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=42);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=42);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=42);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=42);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=42);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111, 22590.10798611111}
TEMP =
  {24.4707, 24.4798, 24.4764, 24.4739, 24.478, 24.4789, 24.4824, 24.4824, 24.4747, 24.4635, 24.4516, 24.4478, 24.4455, 24.4454, 24.4432, 24.4247, 24.4022, 24.3974, 24.3905, 24.3762, 24.3491, 24.3302, 24.3033, 24.2537, 24.2207, 24.2049, 24.176, 24.1546, 24.1347, 24.1181, 24.0707, 23.9718, 23.9707, 23.9759, 23.9664, 23.9393, 23.918, 23.8789, 23.8021, 23.7906, 23.7876, 23.786}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0}
}
