netcdf file-177.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (41 currently)
  variables:
    float LATITUDE(DEPTH=41);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=41);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=41);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=41);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=41);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=41);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926, 22082.25457175926}
TEMP =
  {21.7067, 21.9738, 21.9654, 21.964, 21.9633, 21.9633, 21.9621, 21.9583, 21.9447, 21.935, 21.9135, 21.8938, 21.8761, 21.8235, 21.7288, 21.6726, 21.6294, 21.6164, 21.5892, 21.5819, 21.5675, 21.5542, 21.5286, 21.4934, 21.4464, 21.3828, 21.3268, 21.3062, 21.2801, 21.2502, 21.0053, 20.6918, 20.3995, 20.1796, 20.0168, 19.9424, 19.8366, 19.8069, 19.7806, 19.7359, 19.7238}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0}
}
