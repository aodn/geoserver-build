netcdf file-172.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (28 currently)
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111, 22852.06048611111}
TEMP =
  {21.3355, 21.3195, 21.3203, 21.2978, 21.2823, 21.2767, 21.2732, 21.2573, 21.2439, 21.2365, 21.2324, 21.2293, 21.22, 21.2157, 21.2128, 21.2108, 21.2107, 21.2109, 21.2118, 21.2114, 21.2096, 21.2077, 21.208, 21.2074, 21.2064, 21.2063, 21.2071, 21.2079}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
