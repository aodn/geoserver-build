netcdf file-24.nc {
  dimensions:
    DEPTH = 49;
  variables:
    float LATITUDE(DEPTH=49);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=49);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=49);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=49);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=49);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=49);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556, 22774.143055555556}
TEMP =
  {27.1657, 27.1866, 27.1834, 27.1834, 27.1837, 27.1851, 27.1847, 27.1839, 27.182, 27.1824, 27.1819, 27.1823, 27.1825, 27.1826, 27.1836, 27.1843, 27.1844, 27.185, 27.1865, 27.1865, 27.1866, 27.1856, 27.1839, 27.1828, 27.1832, 27.1832, 27.1837, 27.1841, 27.185, 27.1856, 27.1857, 27.1865, 27.1865, 27.1871, 27.1869, 27.1875, 27.1876, 27.1879, 27.1872, 27.188, 27.1881, 27.1881, 27.1837, 27.1733, 27.1635, 27.1494, 27.1498, 27.1316, 27.1258}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0}
}
