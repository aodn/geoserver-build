netcdf file-156.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518, 22256.053518518518}
TEMP =
  {28.0434, 28.0321, 28.0169, 27.988, 27.8492, 27.5474, 27.3195, 27.1957, 27.155, 27.1396, 27.1324, 27.1297, 27.1286, 27.1276, 27.1264, 27.1257, 27.1249, 27.1245, 27.1241, 27.1238, 27.1239}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853}
}
