netcdf file-151.nc {
  dimensions:
    DEPTH = 23;
  variables:
    float LATITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=23);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=23);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074, 21969.08136574074}
TEMP =
  {29.0324, 28.9632, 28.9349, 28.9204, 28.9096, 28.8969, 28.8849, 28.8736, 28.8679, 28.8666, 28.8656, 28.8645, 28.8632, 28.8619, 28.8604, 28.8585, 28.8562, 28.853, 28.8497, 28.8472, 28.8467, 28.8473, 28.8492}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853}
}
