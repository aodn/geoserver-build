netcdf file-59.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (39 currently)
  variables:
    float LATITUDE(DEPTH=39);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=39);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=39);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=39);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=39);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=39);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416, 115.416}
TIME =
  {23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926, 23147.09832175926}
TEMP =
  {21.1925, 22.0281, 21.7951, 21.7965, 21.7955, 21.7902, 21.7904, 21.7895, 21.7927, 21.7939, 21.7898, 21.7377, 21.7122, 21.6907, 21.6637, 21.5931, 21.4787, 21.309, 21.2242, 21.13, 21.0243, 20.9551, 20.9396, 20.9203, 20.9022, 20.8708, 20.8504, 20.8425, 20.8382, 20.842, 20.8419, 20.832, 20.8251, 20.8192, 20.8161, 20.8145, 20.8131, 20.8125, 20.8183}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0}
}
