netcdf file-25.nc {
  dimensions:
    DEPTH = 47;
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865}
LONGITUDE =
  {113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666}
TIME =
  {22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778, 22884.02215277778}
TEMP =
  {23.8284, 23.8266, 23.8265, 23.8262, 23.8265, 23.8272, 23.8244, 23.8088, 23.7504, 23.6713, 23.6483, 23.6382, 23.6248, 23.6054, 23.5928, 23.5699, 23.5608, 23.5455, 23.5412, 23.5372, 23.5287, 23.534, 23.5323, 23.5264, 23.526, 23.5197, 23.5026, 23.4906, 23.4897, 23.4832, 23.4804, 23.467, 23.4579, 23.4634, 23.4644, 23.4642, 23.471, 23.473, 23.4726, 23.4701, 23.4613, 23.4431, 23.4354, 23.4234, 23.4161, 23.4147, 23.4132}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
