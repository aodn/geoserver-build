netcdf file-43.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (46 currently)
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074, 22517.091261574074}
TEMP =
  {19.8292, 19.829, 19.83, 19.8289, 19.8272, 19.829, 19.8282, 19.8277, 19.8229, 19.8257, 19.8251, 19.8263, 19.8276, 19.8283, 19.8275, 19.8267, 19.8249, 19.8241, 19.8244, 19.8246, 19.8245, 19.8242, 19.8249, 19.8255, 19.8256, 19.8252, 19.8243, 19.8254, 19.8249, 19.8247, 19.8238, 19.8223, 19.8205, 19.811, 19.7948, 19.7951, 19.7824, 19.7633, 19.7367, 19.7163, 19.7083, 19.6991, 19.697, 19.6953, 19.6939, 19.6928}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
