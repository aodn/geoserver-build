netcdf file-126.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (28 currently)
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408, 22944.082094907408}
TEMP =
  {25.4327, 24.9257, 24.9699, 24.9606, 24.9471, 24.9316, 24.9178, 24.911, 24.909, 24.9086, 24.9093, 24.9095, 24.9098, 24.9098, 24.9093, 24.9083, 24.9072, 24.9067, 24.907, 24.9073, 24.9078, 24.9079, 24.9077, 24.9071, 24.9079, 24.9103, 24.9126, 24.9155}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
