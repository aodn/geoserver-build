netcdf IMOS_ANMN-TS_20150113T230000Z_WATR20_FV01_WATR20-1407-Seabird-SBE39-600m-temp-only-150_END-20150122T030000Z_id-7738.nc {
  dimensions:
    TIME = 1177;
  variables:
    double TIME(TIME=1177);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=1177);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=1177);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=1177);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=1177);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=1177);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=1177);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=1177);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=1177);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=1177);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=1177);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=1177);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=1177);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been filled using the DEPTH median (mooring).";
  :instrument = "Seabird         SBE39 [600m] temp only";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "3949303-4138";
  :history = "2015-01-29T06:32:01Z - depthPP: Depth computed from the 2 nearest pressure sensors available, using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 150.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = 0.29053688f; // float
  :geospatial_vertical_max = 161.77881f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-22T03:00:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.965277777777, 23753.972222222223, 23753.979166666668, 23753.98611111111, 23753.993055555555, 23754.0, 23754.006944444445, 23754.01388888889, 23754.020833333332, 23754.027777777777, 23754.034722222223, 23754.041666666668, 23754.04861111111, 23754.055555555555, 23754.0625, 23754.069444444445, 23754.07638888889, 23754.083333333332, 23754.090277777777, 23754.097222222223, 23754.104166666668, 23754.11111111111, 23754.118055555555, 23754.125, 23754.131944444445, 23754.13888888889, 23754.145833333332, 23754.152777777777, 23754.159722222223, 23754.166666666668, 23754.17361111111, 23754.180555555555, 23754.1875, 23754.194444444445, 23754.20138888889, 23754.208333333332, 23754.215277777777, 23754.222222222223, 23754.229166666668, 23754.23611111111, 23754.243055555555, 23754.25, 23754.256944444445, 23754.26388888889, 23754.270833333332, 23754.277777777777, 23754.284722222223, 23754.291666666668, 23754.29861111111, 23754.305555555555, 23754.3125, 23754.319444444445, 23754.32638888889, 23754.333333333332, 23754.340277777777, 23754.347222222223, 23754.354166666668, 23754.36111111111, 23754.368055555555, 23754.375, 23754.381944444445, 23754.38888888889, 23754.395833333332, 23754.402777777777, 23754.409722222223, 23754.416666666668, 23754.42361111111, 23754.430555555555, 23754.4375, 23754.444444444445, 23754.45138888889, 23754.458333333332, 23754.465277777777, 23754.472222222223, 23754.479166666668, 23754.48611111111, 23754.493055555555, 23754.5, 23754.506944444445, 23754.51388888889, 23754.520833333332, 23754.527777777777, 23754.534722222223, 23754.541666666668, 23754.54861111111, 23754.555555555555, 23754.5625, 23754.569444444445, 23754.57638888889, 23754.583333333332, 23754.590277777777, 23754.597222222223, 23754.604166666668, 23754.61111111111, 23754.618055555555, 23754.625, 23754.631944444445, 23754.63888888889, 23754.645833333332, 23754.652777777777, 23754.659722222223, 23754.666666666668, 23754.67361111111, 23754.680555555555, 23754.6875, 23754.694444444445, 23754.70138888889, 23754.708333333332, 23754.715277777777, 23754.722222222223, 23754.729166666668, 23754.73611111111, 23754.743055555555, 23754.75, 23754.756944444445, 23754.76388888889, 23754.770833333332, 23754.777777777777, 23754.784722222223, 23754.791666666668, 23754.79861111111, 23754.805555555555, 23754.8125, 23754.819444444445, 23754.82638888889, 23754.833333333332, 23754.840277777777, 23754.847222222223, 23754.854166666668, 23754.86111111111, 23754.868055555555, 23754.875, 23754.881944444445, 23754.88888888889, 23754.895833333332, 23754.902777777777, 23754.909722222223, 23754.916666666668, 23754.92361111111, 23754.930555555555, 23754.9375, 23754.944444444445, 23754.95138888889, 23754.958333333332, 23754.965277777777, 23754.972222222223, 23754.979166666668, 23754.98611111111, 23754.993055555555, 23755.0, 23755.006944444445, 23755.01388888889, 23755.020833333332, 23755.027777777777, 23755.034722222223, 23755.041666666668, 23755.04861111111, 23755.055555555555, 23755.0625, 23755.069444444445, 23755.07638888889, 23755.083333333332, 23755.090277777777, 23755.097222222223, 23755.104166666668, 23755.11111111111, 23755.118055555555, 23755.125, 23755.131944444445, 23755.13888888889, 23755.145833333332, 23755.152777777777, 23755.159722222223, 23755.166666666668, 23755.17361111111, 23755.180555555555, 23755.1875, 23755.194444444445, 23755.20138888889, 23755.208333333332, 23755.215277777777, 23755.222222222223, 23755.229166666668, 23755.23611111111, 23755.243055555555, 23755.25, 23755.256944444445, 23755.26388888889, 23755.270833333332, 23755.277777777777, 23755.284722222223, 23755.291666666668, 23755.29861111111, 23755.305555555555, 23755.3125, 23755.319444444445, 23755.32638888889, 23755.333333333332, 23755.340277777777, 23755.347222222223, 23755.354166666668, 23755.36111111111, 23755.368055555555, 23755.375, 23755.381944444445, 23755.38888888889, 23755.395833333332, 23755.402777777777, 23755.409722222223, 23755.416666666668, 23755.42361111111, 23755.430555555555, 23755.4375, 23755.444444444445, 23755.45138888889, 23755.458333333332, 23755.465277777777, 23755.472222222223, 23755.479166666668, 23755.48611111111, 23755.493055555555, 23755.5, 23755.506944444445, 23755.51388888889, 23755.520833333332, 23755.527777777777, 23755.534722222223, 23755.541666666668, 23755.54861111111, 23755.555555555555, 23755.5625, 23755.569444444445, 23755.57638888889, 23755.583333333332, 23755.590277777777, 23755.597222222223, 23755.604166666668, 23755.61111111111, 23755.618055555555, 23755.625, 23755.631944444445, 23755.63888888889, 23755.645833333332, 23755.652777777777, 23755.659722222223, 23755.666666666668, 23755.67361111111, 23755.680555555555, 23755.6875, 23755.694444444445, 23755.70138888889, 23755.708333333332, 23755.715277777777, 23755.722222222223, 23755.729166666668, 23755.73611111111, 23755.743055555555, 23755.75, 23755.756944444445, 23755.76388888889, 23755.770833333332, 23755.777777777777, 23755.784722222223, 23755.791666666668, 23755.79861111111, 23755.805555555555, 23755.8125, 23755.819444444445, 23755.82638888889, 23755.833333333332, 23755.840277777777, 23755.847222222223, 23755.854166666668, 23755.86111111111, 23755.868055555555, 23755.875, 23755.881944444445, 23755.88888888889, 23755.895833333332, 23755.902777777777, 23755.909722222223, 23755.916666666668, 23755.92361111111, 23755.930555555555, 23755.9375, 23755.944444444445, 23755.95138888889, 23755.958333333332, 23755.965277777777, 23755.972222222223, 23755.979166666668, 23755.98611111111, 23755.993055555555, 23756.0, 23756.006944444445, 23756.01388888889, 23756.020833333332, 23756.027777777777, 23756.034722222223, 23756.041666666668, 23756.04861111111, 23756.055555555555, 23756.0625, 23756.069444444445, 23756.07638888889, 23756.083333333332, 23756.090277777777, 23756.097222222223, 23756.104166666668, 23756.11111111111, 23756.118055555555, 23756.125, 23756.131944444445, 23756.13888888889, 23756.145833333332, 23756.152777777777, 23756.159722222223, 23756.166666666668, 23756.17361111111, 23756.180555555555, 23756.1875, 23756.194444444445, 23756.20138888889, 23756.208333333332, 23756.215277777777, 23756.222222222223, 23756.229166666668, 23756.23611111111, 23756.243055555555, 23756.25, 23756.256944444445, 23756.26388888889, 23756.270833333332, 23756.277777777777, 23756.284722222223, 23756.291666666668, 23756.29861111111, 23756.305555555555, 23756.3125, 23756.319444444445, 23756.32638888889, 23756.333333333332, 23756.340277777777, 23756.347222222223, 23756.354166666668, 23756.36111111111, 23756.368055555555, 23756.375, 23756.381944444445, 23756.38888888889, 23756.395833333332, 23756.402777777777, 23756.409722222223, 23756.416666666668, 23756.42361111111, 23756.430555555555, 23756.4375, 23756.444444444445, 23756.45138888889, 23756.458333333332, 23756.465277777777, 23756.472222222223, 23756.479166666668, 23756.48611111111, 23756.493055555555, 23756.5, 23756.506944444445, 23756.51388888889, 23756.520833333332, 23756.527777777777, 23756.534722222223, 23756.541666666668, 23756.54861111111, 23756.555555555555, 23756.5625, 23756.569444444445, 23756.57638888889, 23756.583333333332, 23756.590277777777, 23756.597222222223, 23756.604166666668, 23756.61111111111, 23756.618055555555, 23756.625, 23756.631944444445, 23756.63888888889, 23756.645833333332, 23756.652777777777, 23756.659722222223, 23756.666666666668, 23756.67361111111, 23756.680555555555, 23756.6875, 23756.694444444445, 23756.70138888889, 23756.708333333332, 23756.715277777777, 23756.722222222223, 23756.729166666668, 23756.73611111111, 23756.743055555555, 23756.75, 23756.756944444445, 23756.76388888889, 23756.770833333332, 23756.777777777777, 23756.784722222223, 23756.791666666668, 23756.79861111111, 23756.805555555555, 23756.8125, 23756.819444444445, 23756.82638888889, 23756.833333333332, 23756.840277777777, 23756.847222222223, 23756.854166666668, 23756.86111111111, 23756.868055555555, 23756.875, 23756.881944444445, 23756.88888888889, 23756.895833333332, 23756.902777777777, 23756.909722222223, 23756.916666666668, 23756.92361111111, 23756.930555555555, 23756.9375, 23756.944444444445, 23756.95138888889, 23756.958333333332, 23756.965277777777, 23756.972222222223, 23756.979166666668, 23756.98611111111, 23756.993055555555, 23757.0, 23757.006944444445, 23757.01388888889, 23757.020833333332, 23757.027777777777, 23757.034722222223, 23757.041666666668, 23757.04861111111, 23757.055555555555, 23757.0625, 23757.069444444445, 23757.07638888889, 23757.083333333332, 23757.090277777777, 23757.097222222223, 23757.104166666668, 23757.11111111111, 23757.118055555555, 23757.125, 23757.131944444445, 23757.13888888889, 23757.145833333332, 23757.152777777777, 23757.159722222223, 23757.166666666668, 23757.17361111111, 23757.180555555555, 23757.1875, 23757.194444444445, 23757.20138888889, 23757.208333333332, 23757.215277777777, 23757.222222222223, 23757.229166666668, 23757.23611111111, 23757.243055555555, 23757.25, 23757.256944444445, 23757.26388888889, 23757.270833333332, 23757.277777777777, 23757.284722222223, 23757.291666666668, 23757.29861111111, 23757.305555555555, 23757.3125, 23757.319444444445, 23757.32638888889, 23757.333333333332, 23757.340277777777, 23757.347222222223, 23757.354166666668, 23757.36111111111, 23757.368055555555, 23757.375, 23757.381944444445, 23757.38888888889, 23757.395833333332, 23757.402777777777, 23757.409722222223, 23757.416666666668, 23757.42361111111, 23757.430555555555, 23757.4375, 23757.444444444445, 23757.45138888889, 23757.458333333332, 23757.465277777777, 23757.472222222223, 23757.479166666668, 23757.48611111111, 23757.493055555555, 23757.5, 23757.506944444445, 23757.51388888889, 23757.520833333332, 23757.527777777777, 23757.534722222223, 23757.541666666668, 23757.54861111111, 23757.555555555555, 23757.5625, 23757.569444444445, 23757.57638888889, 23757.583333333332, 23757.590277777777, 23757.597222222223, 23757.604166666668, 23757.61111111111, 23757.618055555555, 23757.625, 23757.631944444445, 23757.63888888889, 23757.645833333332, 23757.652777777777, 23757.659722222223, 23757.666666666668, 23757.67361111111, 23757.680555555555, 23757.6875, 23757.694444444445, 23757.70138888889, 23757.708333333332, 23757.715277777777, 23757.722222222223, 23757.729166666668, 23757.73611111111, 23757.743055555555, 23757.75, 23757.756944444445, 23757.76388888889, 23757.770833333332, 23757.777777777777, 23757.784722222223, 23757.791666666668, 23757.79861111111, 23757.805555555555, 23757.8125, 23757.819444444445, 23757.82638888889, 23757.833333333332, 23757.840277777777, 23757.847222222223, 23757.854166666668, 23757.86111111111, 23757.868055555555, 23757.875, 23757.881944444445, 23757.88888888889, 23757.895833333332, 23757.902777777777, 23757.909722222223, 23757.916666666668, 23757.92361111111, 23757.930555555555, 23757.9375, 23757.944444444445, 23757.95138888889, 23757.958333333332, 23757.965277777777, 23757.972222222223, 23757.979166666668, 23757.98611111111, 23757.993055555555, 23758.0, 23758.006944444445, 23758.01388888889, 23758.020833333332, 23758.027777777777, 23758.034722222223, 23758.041666666668, 23758.04861111111, 23758.055555555555, 23758.0625, 23758.069444444445, 23758.07638888889, 23758.083333333332, 23758.090277777777, 23758.097222222223, 23758.104166666668, 23758.11111111111, 23758.118055555555, 23758.125, 23758.131944444445, 23758.13888888889, 23758.145833333332, 23758.152777777777, 23758.159722222223, 23758.166666666668, 23758.17361111111, 23758.180555555555, 23758.1875, 23758.194444444445, 23758.20138888889, 23758.208333333332, 23758.215277777777, 23758.222222222223, 23758.229166666668, 23758.23611111111, 23758.243055555555, 23758.25, 23758.256944444445, 23758.26388888889, 23758.270833333332, 23758.277777777777, 23758.284722222223, 23758.291666666668, 23758.29861111111, 23758.305555555555, 23758.3125, 23758.319444444445, 23758.32638888889, 23758.333333333332, 23758.340277777777, 23758.347222222223, 23758.354166666668, 23758.36111111111, 23758.368055555555, 23758.375, 23758.381944444445, 23758.38888888889, 23758.395833333332, 23758.402777777777, 23758.409722222223, 23758.416666666668, 23758.42361111111, 23758.430555555555, 23758.4375, 23758.444444444445, 23758.45138888889, 23758.458333333332, 23758.465277777777, 23758.472222222223, 23758.479166666668, 23758.48611111111, 23758.493055555555, 23758.5, 23758.506944444445, 23758.51388888889, 23758.520833333332, 23758.527777777777, 23758.534722222223, 23758.541666666668, 23758.54861111111, 23758.555555555555, 23758.5625, 23758.569444444445, 23758.57638888889, 23758.583333333332, 23758.590277777777, 23758.597222222223, 23758.604166666668, 23758.61111111111, 23758.618055555555, 23758.625, 23758.631944444445, 23758.63888888889, 23758.645833333332, 23758.652777777777, 23758.659722222223, 23758.666666666668, 23758.67361111111, 23758.680555555555, 23758.6875, 23758.694444444445, 23758.70138888889, 23758.708333333332, 23758.715277777777, 23758.722222222223, 23758.729166666668, 23758.73611111111, 23758.743055555555, 23758.75, 23758.756944444445, 23758.76388888889, 23758.770833333332, 23758.777777777777, 23758.784722222223, 23758.791666666668, 23758.79861111111, 23758.805555555555, 23758.8125, 23758.819444444445, 23758.82638888889, 23758.833333333332, 23758.840277777777, 23758.847222222223, 23758.854166666668, 23758.86111111111, 23758.868055555555, 23758.875, 23758.881944444445, 23758.88888888889, 23758.895833333332, 23758.902777777777, 23758.909722222223, 23758.916666666668, 23758.92361111111, 23758.930555555555, 23758.9375, 23758.944444444445, 23758.95138888889, 23758.958333333332, 23758.965277777777, 23758.972222222223, 23758.979166666668, 23758.98611111111, 23758.993055555555, 23759.0, 23759.006944444445, 23759.01388888889, 23759.020833333332, 23759.027777777777, 23759.034722222223, 23759.041666666668, 23759.04861111111, 23759.055555555555, 23759.0625, 23759.069444444445, 23759.07638888889, 23759.083333333332, 23759.090277777777, 23759.097222222223, 23759.104166666668, 23759.11111111111, 23759.118055555555, 23759.125, 23759.131944444445, 23759.13888888889, 23759.145833333332, 23759.152777777777, 23759.159722222223, 23759.166666666668, 23759.17361111111, 23759.180555555555, 23759.1875, 23759.194444444445, 23759.20138888889, 23759.208333333332, 23759.215277777777, 23759.222222222223, 23759.229166666668, 23759.23611111111, 23759.243055555555, 23759.25, 23759.256944444445, 23759.26388888889, 23759.270833333332, 23759.277777777777, 23759.284722222223, 23759.291666666668, 23759.29861111111, 23759.305555555555, 23759.3125, 23759.319444444445, 23759.32638888889, 23759.333333333332, 23759.340277777777, 23759.347222222223, 23759.354166666668, 23759.36111111111, 23759.368055555555, 23759.375, 23759.381944444445, 23759.38888888889, 23759.395833333332, 23759.402777777777, 23759.409722222223, 23759.416666666668, 23759.42361111111, 23759.430555555555, 23759.4375, 23759.444444444445, 23759.45138888889, 23759.458333333332, 23759.465277777777, 23759.472222222223, 23759.479166666668, 23759.48611111111, 23759.493055555555, 23759.5, 23759.506944444445, 23759.51388888889, 23759.520833333332, 23759.527777777777, 23759.534722222223, 23759.541666666668, 23759.54861111111, 23759.555555555555, 23759.5625, 23759.569444444445, 23759.57638888889, 23759.583333333332, 23759.590277777777, 23759.597222222223, 23759.604166666668, 23759.61111111111, 23759.618055555555, 23759.625, 23759.631944444445, 23759.63888888889, 23759.645833333332, 23759.652777777777, 23759.659722222223, 23759.666666666668, 23759.67361111111, 23759.680555555555, 23759.6875, 23759.694444444445, 23759.70138888889, 23759.708333333332, 23759.715277777777, 23759.722222222223, 23759.729166666668, 23759.73611111111, 23759.743055555555, 23759.75, 23759.756944444445, 23759.76388888889, 23759.770833333332, 23759.777777777777, 23759.784722222223, 23759.791666666668, 23759.79861111111, 23759.805555555555, 23759.8125, 23759.819444444445, 23759.82638888889, 23759.833333333332, 23759.840277777777, 23759.847222222223, 23759.854166666668, 23759.86111111111, 23759.868055555555, 23759.875, 23759.881944444445, 23759.88888888889, 23759.895833333332, 23759.902777777777, 23759.909722222223, 23759.916666666668, 23759.92361111111, 23759.930555555555, 23759.9375, 23759.944444444445, 23759.95138888889, 23759.958333333332, 23759.965277777777, 23759.972222222223, 23759.979166666668, 23759.98611111111, 23759.993055555555, 23760.0, 23760.006944444445, 23760.01388888889, 23760.020833333332, 23760.027777777777, 23760.034722222223, 23760.041666666668, 23760.04861111111, 23760.055555555555, 23760.0625, 23760.069444444445, 23760.07638888889, 23760.083333333332, 23760.090277777777, 23760.097222222223, 23760.104166666668, 23760.11111111111, 23760.118055555555, 23760.125, 23760.131944444445, 23760.13888888889, 23760.145833333332, 23760.152777777777, 23760.159722222223, 23760.166666666668, 23760.17361111111, 23760.180555555555, 23760.1875, 23760.194444444445, 23760.20138888889, 23760.208333333332, 23760.215277777777, 23760.222222222223, 23760.229166666668, 23760.23611111111, 23760.243055555555, 23760.25, 23760.256944444445, 23760.26388888889, 23760.270833333332, 23760.277777777777, 23760.284722222223, 23760.291666666668, 23760.29861111111, 23760.305555555555, 23760.3125, 23760.319444444445, 23760.32638888889, 23760.333333333332, 23760.340277777777, 23760.347222222223, 23760.354166666668, 23760.36111111111, 23760.368055555555, 23760.375, 23760.381944444445, 23760.38888888889, 23760.395833333332, 23760.402777777777, 23760.409722222223, 23760.416666666668, 23760.42361111111, 23760.430555555555, 23760.4375, 23760.444444444445, 23760.45138888889, 23760.458333333332, 23760.465277777777, 23760.472222222223, 23760.479166666668, 23760.48611111111, 23760.493055555555, 23760.5, 23760.506944444445, 23760.51388888889, 23760.520833333332, 23760.527777777777, 23760.534722222223, 23760.541666666668, 23760.54861111111, 23760.555555555555, 23760.5625, 23760.569444444445, 23760.57638888889, 23760.583333333332, 23760.590277777777, 23760.597222222223, 23760.604166666668, 23760.61111111111, 23760.618055555555, 23760.625, 23760.631944444445, 23760.63888888889, 23760.645833333332, 23760.652777777777, 23760.659722222223, 23760.666666666668, 23760.67361111111, 23760.680555555555, 23760.6875, 23760.694444444445, 23760.70138888889, 23760.708333333332, 23760.715277777777, 23760.722222222223, 23760.729166666668, 23760.73611111111, 23760.743055555555, 23760.75, 23760.756944444445, 23760.76388888889, 23760.770833333332, 23760.777777777777, 23760.784722222223, 23760.791666666668, 23760.79861111111, 23760.805555555555, 23760.8125, 23760.819444444445, 23760.82638888889, 23760.833333333332, 23760.840277777777, 23760.847222222223, 23760.854166666668, 23760.86111111111, 23760.868055555555, 23760.875, 23760.881944444445, 23760.88888888889, 23760.895833333332, 23760.902777777777, 23760.909722222223, 23760.916666666668, 23760.92361111111, 23760.930555555555, 23760.9375, 23760.944444444445, 23760.95138888889, 23760.958333333332, 23760.965277777777, 23760.972222222223, 23760.979166666668, 23760.98611111111, 23760.993055555555, 23761.0, 23761.006944444445, 23761.01388888889, 23761.020833333332, 23761.027777777777, 23761.034722222223, 23761.041666666668, 23761.04861111111, 23761.055555555555, 23761.0625, 23761.069444444445, 23761.07638888889, 23761.083333333332, 23761.090277777777, 23761.097222222223, 23761.104166666668, 23761.11111111111, 23761.118055555555, 23761.125, 23761.131944444445, 23761.13888888889, 23761.145833333332, 23761.152777777777, 23761.159722222223, 23761.166666666668, 23761.17361111111, 23761.180555555555, 23761.1875, 23761.194444444445, 23761.20138888889, 23761.208333333332, 23761.215277777777, 23761.222222222223, 23761.229166666668, 23761.23611111111, 23761.243055555555, 23761.25, 23761.256944444445, 23761.26388888889, 23761.270833333332, 23761.277777777777, 23761.284722222223, 23761.291666666668, 23761.29861111111, 23761.305555555555, 23761.3125, 23761.319444444445, 23761.32638888889, 23761.333333333332, 23761.340277777777, 23761.347222222223, 23761.354166666668, 23761.36111111111, 23761.368055555555, 23761.375, 23761.381944444445, 23761.38888888889, 23761.395833333332, 23761.402777777777, 23761.409722222223, 23761.416666666668, 23761.42361111111, 23761.430555555555, 23761.4375, 23761.444444444445, 23761.45138888889, 23761.458333333332, 23761.465277777777, 23761.472222222223, 23761.479166666668, 23761.48611111111, 23761.493055555555, 23761.5, 23761.506944444445, 23761.51388888889, 23761.520833333332, 23761.527777777777, 23761.534722222223, 23761.541666666668, 23761.54861111111, 23761.555555555555, 23761.5625, 23761.569444444445, 23761.57638888889, 23761.583333333332, 23761.590277777777, 23761.597222222223, 23761.604166666668, 23761.61111111111, 23761.618055555555, 23761.625, 23761.631944444445, 23761.63888888889, 23761.645833333332, 23761.652777777777, 23761.659722222223, 23761.666666666668, 23761.67361111111, 23761.680555555555, 23761.6875, 23761.694444444445, 23761.70138888889, 23761.708333333332, 23761.715277777777, 23761.722222222223, 23761.729166666668, 23761.73611111111, 23761.743055555555, 23761.75, 23761.756944444445, 23761.76388888889, 23761.770833333332, 23761.777777777777, 23761.784722222223, 23761.791666666668, 23761.79861111111, 23761.805555555555, 23761.8125, 23761.819444444445, 23761.82638888889, 23761.833333333332, 23761.840277777777, 23761.847222222223, 23761.854166666668, 23761.86111111111, 23761.868055555555, 23761.875, 23761.881944444445, 23761.88888888889, 23761.895833333332, 23761.902777777777, 23761.909722222223, 23761.916666666668, 23761.92361111111, 23761.930555555555, 23761.9375, 23761.944444444445, 23761.95138888889, 23761.958333333332, 23761.965277777777, 23761.972222222223, 23761.979166666668, 23761.98611111111, 23761.993055555555, 23762.0, 23762.006944444445, 23762.01388888889, 23762.020833333332, 23762.027777777777, 23762.034722222223, 23762.041666666668, 23762.04861111111, 23762.055555555555, 23762.0625, 23762.069444444445, 23762.07638888889, 23762.083333333332, 23762.090277777777, 23762.097222222223, 23762.104166666668, 23762.11111111111, 23762.118055555555, 23762.125}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =150.0
TEMP =
  {16.8141, 16.886, 16.9306, 16.9891, 16.9635, 16.9696, 16.9278, 16.919, 16.9169, 16.8956, 17.0687, 17.1063, 16.9637, 16.991, 17.0828, 17.1216, 17.071, 17.1688, 17.1157, 17.1407, 17.1623, 17.1892, 17.2314, 17.2401, 17.2426, 17.2622, 17.2831, 17.2285, 17.1767, 17.1963, 17.1678, 17.2072, 17.2445, 17.2028, 17.1604, 17.1354, 17.1523, 17.1446, 17.1379, 17.1347, 17.1355, 17.1292, 17.1292, 17.1426, 17.136, 17.157, 17.1463, 17.2133, 17.1857, 17.0781, 17.1119, 17.118, 17.1309, 17.1779, 17.0842, 17.1146, 17.1516, 17.2421, 17.2208, 17.1434, 17.1258, 17.1775, 17.086, 17.0863, 17.0801, 17.0608, 17.02, 17.0447, 17.2096, 17.1787, 17.1987, 17.2115, 17.1664, 17.1111, 17.1075, 17.0981, 17.1863, 17.3269, 17.3264, 17.3165, 17.2666, 17.2863, 17.3626, 17.2506, 17.2655, 17.2564, 17.4303, 17.4506, 17.2627, 17.1684, 17.156, 17.4623, 17.1047, 17.0496, 17.0753, 17.0871, 17.4538, 17.3945, 17.3629, 17.3409, 17.3333, 17.3228, 17.279, 17.308, 17.3396, 17.338, 17.4418, 17.4209, 17.4414, 17.5888, 17.7173, 17.7115, 17.6641, 17.4592, 17.4327, 17.4191, 17.393, 17.3294, 17.3127, 17.4297, 17.4335, 17.4249, 17.4797, 17.4765, 17.4611, 17.4496, 17.4303, 17.4225, 17.4159, 17.4019, 17.4073, 17.4008, 17.3816, 17.3663, 17.3789, 17.3684, 17.3241, 17.3126, 17.3332, 17.3207, 17.3084, 17.3431, 17.3508, 17.3511, 17.35, 17.3423, 17.2956, 17.2746, 17.2699, 17.267, 17.2946, 17.3604, 17.4667, 17.5111, 17.5006, 17.5147, 17.519, 17.5957, 17.6777, 17.6771, 17.67, 17.6234, 17.6841, 17.5914, 17.5667, 17.5796, 17.5803, 17.5038, 17.5106, 17.6075, 17.7187, 17.6749, 17.6393, 17.7987, 17.8384, 17.8453, 17.8643, 17.8392, 17.7502, 17.5687, 17.5378, 17.5216, 17.5681, 17.5872, 17.6265, 17.6837, 17.7216, 17.7199, 17.7368, 17.8439, 17.8179, 17.8582, 17.849, 17.8539, 17.7665, 17.7299, 17.7329, 17.7556, 17.7512, 17.7735, 17.8539, 17.8621, 17.8651, 17.8613, 17.8612, 17.8285, 17.8487, 17.8567, 17.8345, 17.8733, 17.8893, 17.8716, 17.881, 17.7872, 17.836, 17.913, 17.8958, 17.9163, 17.9102, 17.9023, 17.8658, 17.7867, 17.7923, 17.8921, 17.9052, 17.9412, 17.8994, 17.8857, 17.8955, 17.8969, 17.8953, 17.8955, 17.9009, 17.8875, 17.8856, 17.9355, 17.8937, 17.9091, 17.8784, 17.8745, 17.8884, 17.8707, 17.8812, 17.8774, 17.8717, 17.8848, 17.8841, 17.9026, 17.9039, 17.9579, 17.976, 17.9911, 17.9874, 17.9699, 17.9704, 17.9587, 17.9321, 17.9294, 17.9627, 17.9677, 17.9637, 17.981, 17.9794, 17.9753, 17.9453, 17.9068, 17.9355, 17.9603, 17.9503, 17.9361, 17.8841, 17.823, 17.8082, 17.7414, 17.6486, 17.6169, 17.5633, 17.5926, 17.5938, 17.5646, 17.6262, 17.6873, 17.768, 17.8334, 17.858, 17.6455, 17.5282, 17.5048, 17.4986, 17.5141, 17.5215, 17.6331, 17.4976, 17.4834, 17.6526, 17.5711, 17.5275, 17.707, 17.7348, 17.5332, 17.5276, 17.4849, 17.4607, 17.4353, 17.4779, 17.4713, 17.6063, 17.5996, 17.7217, 17.7901, 17.8052, 17.8396, 17.8536, 17.8797, 17.9108, 17.9495, 18.0323, 18.1842, 18.2044, 18.1737, 18.1935, 18.1996, 18.1931, 18.1542, 18.0076, 17.8834, 17.8925, 17.8675, 17.8812, 17.8595, 17.8595, 17.8569, 17.8551, 17.8513, 17.8488, 17.8175, 17.8133, 17.8157, 17.8248, 17.8417, 17.8501, 17.8498, 17.8485, 17.7919, 17.7167, 17.7115, 17.7139, 17.6853, 17.5958, 17.6122, 17.6538, 17.6672, 17.7195, 17.8007, 17.8141, 17.7661, 17.5948, 17.7071, 17.5077, 17.4721, 17.5374, 17.4659, 17.5153, 17.4716, 17.4585, 17.3136, 17.4127, 17.5818, 17.4977, 17.4446, 17.5612, 17.4279, 17.5206, 17.5576, 17.581, 17.5744, 17.5734, 17.5796, 17.5871, 17.7285, 17.7455, 17.7424, 17.7474, 17.7541, 17.7445, 17.7443, 17.653, 17.5846, 17.5805, 17.5916, 17.59, 17.5438, 17.5562, 17.5627, 17.5604, 17.5477, 17.5536, 17.5875, 17.5573, 17.5136, 17.467, 17.5923, 17.6105, 17.7046, 17.6195, 17.6932, 17.6216, 17.5671, 17.5571, 17.5386, 17.6537, 17.6825, 17.6777, 17.5814, 17.5872, 17.5951, 17.6795, 17.6945, 17.6171, 17.6543, 17.6733, 17.6757, 17.5758, 17.5306, 17.4667, 17.4509, 17.4227, 17.4973, 17.4788, 17.3553, 16.8862, 17.1947, 16.7875, 17.0198, 17.2466, 17.2537, 17.2366, 16.9744, 16.5518, 17.0388, 17.0968, 16.9073, 17.1765, 17.3081, 17.2272, 16.9364, 16.818, 16.6687, 17.107, 17.2136, 17.2464, 17.337, 17.4752, 17.4478, 17.4852, 17.4659, 17.4475, 17.4358, 17.4481, 17.3681, 17.4001, 17.455, 17.4255, 17.4156, 17.4878, 17.4438, 17.4483, 17.3675, 17.3304, 17.5075, 17.4936, 17.6871, 17.7136, 17.7152, 17.7167, 17.6205, 17.7064, 17.7383, 17.7516, 17.7619, 17.4455, 17.5068, 17.5586, 17.5632, 17.6853, 17.6725, 17.5003, 17.4801, 17.3947, 17.3582, 17.7301, 17.462, 17.5703, 17.6111, 17.6002, 17.5441, 17.3982, 17.1212, 17.129, 17.0846, 17.068, 16.7101, 17.026, 17.0239, 17.0156, 16.6941, 15.9576, 15.7793, 15.8348, 15.8717, 16.0625, 16.1155, 16.2641, 16.3998, 16.3441, 16.3469, 16.2325, 16.3299, 16.2903, 15.99, 16.0034, 16.2172, 16.2263, 16.0554, 16.1395, 16.131, 16.2204, 16.2774, 16.3364, 16.3305, 16.2756, 16.2394, 16.2332, 16.3612, 16.5646, 16.6321, 16.7031, 16.4552, 16.3914, 16.3556, 16.4593, 16.4182, 16.3647, 16.4609, 16.5337, 16.5658, 16.7209, 16.7081, 16.7158, 16.5816, 16.6503, 16.6921, 16.7264, 16.6811, 16.695, 16.5863, 16.6736, 16.5577, 16.5368, 16.531, 16.5339, 16.7546, 16.7462, 16.7271, 16.5196, 16.4928, 16.4867, 16.481, 16.4766, 16.4666, 16.4583, 16.503, 16.7629, 16.4923, 16.4198, 16.4311, 16.4179, 16.4646, 16.6769, 16.4788, 16.4155, 16.3331, 16.4, 16.4305, 16.4132, 16.3277, 16.2303, 15.9736, 15.9791, 16.0493, 16.1615, 16.1915, 16.1614, 16.1565, 16.3165, 16.3643, 16.3803, 16.3808, 16.3519, 16.2918, 16.3265, 16.3307, 16.3307, 16.3208, 16.3004, 16.319, 16.3255, 16.3235, 16.3315, 16.3169, 16.3665, 16.3997, 16.571, 16.9472, 16.956, 16.948, 16.9496, 17.0006, 17.0192, 17.1052, 17.0111, 16.9807, 16.9371, 16.9691, 16.9848, 16.9968, 16.9552, 16.9415, 16.9203, 16.898, 16.7364, 16.6967, 16.7347, 16.7961, 16.7282, 16.4403, 16.429, 16.5331, 16.6861, 16.6068, 16.4717, 16.6618, 16.6826, 16.6521, 16.5989, 16.3682, 16.3644, 16.3847, 16.3587, 16.2448, 16.2977, 16.2986, 16.2817, 16.2604, 16.2535, 16.2335, 16.2089, 16.1772, 16.2161, 16.2026, 16.2115, 16.2058, 16.243, 16.2773, 16.1566, 16.1783, 16.1515, 16.1332, 16.1794, 16.1811, 16.1734, 16.1664, 16.1545, 16.1482, 16.1272, 16.1213, 16.1077, 16.0962, 16.1149, 16.0811, 16.0507, 16.067, 16.0848, 16.0967, 16.0835, 16.0957, 16.1053, 16.1157, 16.1159, 16.1273, 16.1388, 16.1688, 16.2843, 16.7537, 16.7061, 16.6372, 16.7539, 16.7831, 16.4784, 16.3946, 16.3473, 16.1822, 16.153, 16.1606, 16.1573, 16.1404, 16.1684, 16.1922, 16.3854, 16.4649, 16.4836, 16.6079, 16.5887, 16.578, 16.5851, 16.5434, 16.7811, 16.6396, 16.8046, 16.8244, 16.8225, 16.8254, 16.8157, 16.8184, 16.8342, 16.9147, 16.9383, 17.0241, 17.0586, 16.9792, 16.9266, 16.9652, 16.9949, 16.9253, 16.9817, 17.2024, 17.2585, 17.2015, 17.0644, 17.1096, 17.1391, 17.1057, 17.0657, 17.1015, 17.1005, 17.1313, 17.3695, 17.4219, 17.4146, 17.4115, 17.4053, 17.4716, 17.56, 17.6314, 17.6324, 17.6287, 17.6209, 17.6078, 17.5729, 17.5047, 17.3785, 17.3226, 17.5522, 17.584, 17.5255, 16.9009, 17.3187, 17.3398, 16.997, 17.5087, 17.3309, 17.4947, 17.4969, 17.5183, 17.5382, 17.5433, 17.4039, 17.396, 17.5313, 17.3549, 17.2928, 17.3407, 17.3444, 17.4193, 17.3845, 17.3738, 17.4254, 17.4274, 17.4057, 17.3822, 17.4174, 17.515, 17.5259, 17.4843, 17.4075, 17.4438, 17.456, 17.3566, 17.429, 17.5186, 17.5024, 17.4938, 17.6836, 17.2916, 17.1248, 17.147, 17.0277, 17.1805, 17.1984, 16.9896, 17.2759, 17.624, 17.3894, 17.24, 17.0759, 16.6687, 17.1584, 17.1666, 17.3339, 17.3402, 17.3663, 17.2964, 17.3139, 17.2772, 17.0508, 17.0008, 16.909, 17.0455, 17.1679, 17.1068, 17.0491, 16.6456, 16.9039, 17.0108, 16.739, 16.6643, 16.6508, 16.9933, 17.014, 16.7717, 16.4847, 16.9051, 16.9589, 17.1007, 16.9031, 16.6526, 16.5397, 16.6314, 16.7234, 16.6602, 16.1352, 16.5222, 16.3192, 16.9126, 16.5322, 17.2025, 16.3165, 16.3042, 16.3745, 16.2218, 16.254, 16.2909, 16.8471, 16.6922, 17.0039, 16.987, 16.95, 16.6852, 16.2374, 16.2643, 16.7556, 16.4053, 16.9286, 17.3636, 16.8734, 17.3597, 17.4559, 17.4346, 17.4483, 17.4359, 17.335, 17.2284, 17.2196, 17.1772, 17.1166, 17.094, 17.0941, 21.2863, 23.1813, 25.6225, 24.2833, 23.7603, 23.6397, 23.8418, 22.7021, 22.3071, 22.2357, 22.39, 22.2589, 22.2498, 22.2063, 22.1865, 22.5211, 23.5603, 24.9208, 26.3503, 28.0559, 28.0342, 27.959, 27.9421, 27.8298, 27.8228, 27.8037, 27.7752, 27.7446, 27.7092, 27.6704, 27.6259, 27.5716, 27.5118, 27.447, 27.3777, 27.3046, 27.2311, 27.1572, 27.0857, 27.0134, 26.9406, 26.8627, 26.7868, 26.7106, 26.635, 26.5624, 26.4905, 26.4205, 26.3517, 26.2819, 26.2102, 26.1373, 26.0661, 25.9892, 25.9109, 25.8297, 25.7465, 25.6644, 25.5841, 25.5055, 25.4291, 25.3533, 25.2783, 25.2055, 25.1346, 25.0658, 24.9998, 24.9347, 24.8728, 24.8106, 24.7535, 24.6935, 24.6364, 24.5785, 24.5213, 24.4651, 24.4054, 24.3432, 24.2794, 24.2137, 24.1452, 24.0715, 23.9952, 23.9205, 23.8471, 23.7798, 23.7191, 23.6662, 23.6157, 23.5684, 23.5258, 23.4829, 23.4368, 23.3875, 23.3342, 23.2802, 23.2257, 23.169, 23.1113, 23.055, 22.9979, 22.9397, 22.8795, 22.8193, 22.7602, 22.7024, 22.6446, 22.5885, 22.532, 22.4765, 22.4206, 22.3647, 22.3084, 22.2521, 22.1955, 22.139, 22.0832, 22.0293, 21.9782, 21.9279, 21.8807, 21.8353, 21.7923, 21.7493, 21.7091, 21.6725, 21.636, 21.6037, 21.573, 21.5438, 21.5141, 21.4881, 21.4619, 21.4399, 21.422, 21.4076, 21.3965, 21.3877, 21.3811, 21.3761, 21.3731, 21.3723, 21.3715, 21.3719, 21.3755, 21.3787, 21.3862, 21.3944, 21.4048, 21.4197, 21.4534, 21.6424, 21.8574, 22.0134, 22.2791, 22.3167, 22.6532, 22.9016, 23.048, 23.6872, 24.0412, 24.3173, 24.518, 24.723, 25.1683, 25.4446, 25.6101, 25.7547, 25.8619, 25.9551, 25.9606, 25.7794, 25.5817, 25.4161, 25.2686, 25.1385, 25.0232, 24.9213, 24.83, 24.7478, 24.6758, 24.6101, 24.5676, 24.539, 24.5155, 24.4974, 24.483, 24.4732, 24.4666, 24.462, 24.4592, 24.459, 24.4612, 24.4641, 24.4679, 24.472, 24.4767, 24.4812, 24.4859, 24.4918, 24.4969, 24.502, 24.5083, 24.5123, 24.5167, 24.523, 24.5272, 24.531, 24.5372, 24.5417, 24.5459, 24.5504, 24.5541, 24.5584, 24.5627, 24.5666, 24.5706, 24.5754, 24.5791, 24.5833, 24.5869, 24.5914, 24.5952, 24.5992, 24.6037, 24.6077, 24.6119, 24.6152, 24.6188, 24.6222, 24.6259, 24.6286, 24.6315, 24.6353, 24.6368, 24.6396, 24.642, 24.6436, 24.6464, 24.6475, 24.6509, 24.6519, 24.6531, 24.6542, 24.656, 24.6574, 24.6585, 24.6586, 24.6604, 24.662, 24.6624, 24.6631, 24.6642, 24.6645, 24.6664, 24.6383, 24.617, 24.5983, 24.5771, 24.5502, 24.5253, 24.5045, 24.4867, 24.4687, 24.4494, 24.4269, 24.4055, 24.3885, 24.3748, 24.3624, 24.3489, 24.3235, 24.3057, 24.2859, 24.2656, 24.246, 24.2289, 24.2137, 24.1992, 24.182, 24.1719, 24.1598, 24.1461, 24.1364, 24.1295, 24.1201, 24.1149, 24.1057, 24.0999, 24.0877}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_REL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
DEPTH =
  {161.27293, 161.17195, 161.18497, 161.19687, 161.23277, 161.20917, 161.20578, 161.21088, 161.18484, 161.20737, 161.28072, 161.21616, 161.21121, 161.28601, 161.20724, 161.29405, 161.26804, 161.21977, 161.30804, 161.29651, 161.23839, 161.33878, 161.32346, 161.34549, 161.35637, 161.36447, 161.33516, 161.28622, 161.33675, 161.31384, 161.32687, 161.30666, 161.34781, 161.36935, 161.39365, 161.387, 161.4149, 161.41844, 161.3981, 161.40399, 161.39774, 161.45035, 161.43085, 161.37257, 161.44897, 161.40399, 161.4226, 161.41214, 161.44386, 161.3963, 161.46445, 161.46387, 161.47821, 161.50089, 161.45087, 161.48196, 161.43619, 161.40869, 161.48007, 161.47537, 161.44315, 161.44878, 161.50964, 161.48135, 161.46109, 161.5135, 161.45514, 161.46025, 161.46648, 161.45697, 161.48463, 161.47089, 161.48346, 161.50903, 161.48123, 161.49773, 161.48882, 161.40094, 161.47723, 161.44424, 161.41377, 161.40018, 161.45529, 161.43791, 161.3716, 161.43799, 161.36325, 161.39253, 161.36841, 161.38086, 161.35155, 161.37328, 161.38084, 161.36568, 161.37842, 161.33133, 161.28986, 161.30089, 161.27461, 161.25377, 161.25256, 161.25136, 161.28967, 161.2192, 161.19077, 161.29291, 161.21957, 161.25339, 161.21243, 161.22037, 161.23672, 161.26144, 161.26869, 161.21373, 161.20494, 161.1885, 161.19095, 161.15024, 161.14572, 161.16318, 161.15369, 161.15742, 161.1347, 161.15091, 161.09924, 161.13303, 161.10123, 161.14597, 161.15701, 161.07693, 161.15388, 161.08972, 161.15918, 161.1309, 161.07245, 161.0698, 161.08426, 161.053, 161.12497, 161.11076, 161.06612, 161.12576, 161.09436, 161.11855, 161.1295, 161.14102, 161.09969, 161.14006, 161.11801, 161.17152, 161.20319, 161.16907, 161.16779, 161.1601, 161.18889, 161.15045, 161.18655, 161.19287, 161.2066, 161.20384, 161.23431, 161.23618, 161.27379, 161.22913, 161.259, 161.21109, 161.25647, 161.26985, 161.31181, 161.24312, 161.26251, 161.28094, 161.28818, 161.30405, 161.25943, 161.3211, 161.29588, 161.26093, 161.26437, 161.30832, 161.38937, 161.3474, 161.34195, 161.39703, 161.35101, 161.3328, 161.3748, 161.40161, 161.35864, 161.3686, 161.3368, 161.40964, 161.43842, 161.39258, 161.40262, 161.44017, 161.4234, 161.4216, 161.47058, 161.45328, 161.48663, 161.44559, 161.43494, 161.50162, 161.48709, 161.4807, 161.46042, 161.45358, 161.49571, 161.50906, 161.496, 161.4536, 161.49615, 161.51312, 161.45914, 161.48389, 161.44812, 161.51343, 161.44473, 161.46933, 161.46886, 161.45221, 161.40271, 161.413, 161.41527, 161.4166, 161.38742, 161.42538, 161.4198, 161.37347, 161.37427, 161.32819, 161.42268, 161.29645, 161.36841, 161.34384, 161.30536, 161.31137, 161.29724, 161.28383, 161.25327, 161.23727, 161.20065, 161.24335, 161.22208, 161.16788, 161.16309, 161.1659, 161.17914, 161.14207, 161.23303, 161.15396, 161.10217, 161.11096, 161.18903, 161.13614, 161.04477, 161.08432, 161.14407, 161.08398, 161.1238, 161.08034, 161.11014, 161.03592, 161.05997, 161.03365, 161.04398, 161.06715, 161.04541, 161.05731, 161.03842, 161.09677, 161.07632, 161.08173, 161.06314, 161.10599, 161.0591, 161.13771, 161.05118, 161.00998, 161.09918, 161.09781, 161.11627, 161.07164, 161.1075, 161.10727, 161.09897, 161.12578, 161.1341, 161.1901, 161.11594, 161.132, 161.14838, 161.18167, 161.15921, 161.16376, 161.19756, 161.16875, 161.18835, 161.24588, 161.20792, 161.17824, 161.22148, 161.27115, 161.27893, 161.24493, 161.24908, 161.30551, 161.27576, 161.26569, 161.27014, 161.32298, 161.25381, 161.1856, 161.27936, 161.3114, 161.31882, 161.28326, 161.32388, 161.29532, 161.28865, 161.37659, 161.36267, 161.27249, 161.34454, 161.35211, 161.3067, 161.37523, 161.36761, 161.3255, 161.39926, 161.4017, 161.38712, 161.44016, 161.42764, 161.39957, 161.43584, 161.42384, 161.47144, 161.47144, 161.51962, 161.48764, 161.53615, 161.51393, 161.51976, 161.49292, 161.55682, 161.56348, 161.56976, 161.57974, 161.538, 161.58746, 161.5682, 161.6062, 161.51938, 161.57303, 161.58432, 161.57906, 161.54176, 161.54453, 161.56128, 161.61343, 161.58824, 161.62123, 161.63116, 161.5087, 161.52179, 161.52704, 161.6061, 161.51723, 161.49611, 161.5203, 161.52054, 161.48128, 161.49786, 161.47516, 161.54503, 161.491, 161.40561, 161.4299, 161.41083, 161.37799, 161.35004, 161.3676, 161.30435, 161.34818, 161.31345, 161.33218, 161.26132, 161.27388, 161.24965, 161.25858, 161.16487, 161.24472, 161.20122, 161.16437, 161.16545, 161.16798, 161.1939, 161.14542, 161.11874, 161.15369, 161.05116, 161.10226, 161.09747, 161.03506, 160.99258, 161.10825, 161.08432, 161.0459, 160.9982, 161.09982, 160.99695, 161.0047, 161.0854, 161.12123, 161.09155, 161.05809, 161.00946, 161.09134, 161.08215, 161.03796, 161.02502, 161.08269, 161.04037, 161.06189, 161.1141, 161.06427, 161.108, 161.08344, 161.09065, 161.03604, 161.07547, 161.1333, 161.10608, 161.12128, 161.14386, 161.12717, 161.11984, 161.11928, 161.13371, 161.21558, 161.2058, 161.1694, 161.21977, 161.22995, 161.19908, 161.23572, 161.2437, 161.24493, 161.28607, 161.24716, 161.29453, 161.27571, 161.258, 161.31586, 161.29446, 161.29066, 161.318, 161.36804, 161.29941, 161.34813, 161.32018, 161.38275, 161.27667, 161.38658, 161.30809, 161.37323, 161.34537, 161.36523, 161.34274, 161.3375, 161.39145, 161.39877, 161.47018, 161.44803, 161.4088, 161.42163, 161.44637, 161.4131, 161.46478, 161.43799, 161.52481, 161.55275, 161.5069, 161.52365, 161.56494, 161.62517, 161.59508, 161.52579, 161.53639, 161.59175, 161.64784, 161.63933, 161.63686, 161.58092, 161.60567, 161.67206, 161.65971, 161.74242, 161.66095, 161.66994, 161.75235, 161.6725, 161.65642, 161.72623, 161.73825, 161.66116, 161.68863, 161.63608, 161.69028, 161.68259, 161.65738, 161.63991, 161.67606, 161.63145, 161.58344, 161.58904, 161.65138, 161.56422, 161.61989, 161.62503, 161.53513, 161.56451, 161.52075, 161.45107, 161.47595, 161.51224, 161.38339, 161.40689, 161.39505, 161.3381, 161.36713, 161.32828, 161.33234, 161.294, 161.30328, 161.27548, 161.23227, 161.27776, 161.22607, 161.22455, 161.14969, 161.15268, 161.08815, 161.18576, 161.06906, 161.09488, 161.06284, 161.0991, 161.052, 160.98053, 161.05292, 161.14575, 161.05995, 160.9907, 161.0712, 161.02042, 161.05716, 161.02339, 161.01318, 161.05635, 160.96907, 161.02138, 161.09076, 160.98566, 161.05048, 161.07484, 161.00757, 161.0788, 161.09485, 161.08264, 161.10498, 161.01404, 161.02309, 161.05948, 161.10278, 161.12868, 161.09755, 161.1334, 161.16904, 161.18927, 161.17482, 161.17181, 161.18028, 161.16205, 161.20267, 161.2524, 161.26355, 161.29968, 161.31519, 161.298, 161.31754, 161.26976, 161.24991, 161.30603, 161.33083, 161.25853, 161.32124, 161.38062, 161.30652, 161.34384, 161.28688, 161.35098, 161.3003, 161.32639, 161.26868, 161.33694, 161.36191, 161.3744, 161.32462, 161.34644, 161.35669, 161.34283, 161.40643, 161.45224, 161.48965, 161.41022, 161.45935, 161.42517, 161.44647, 161.44008, 161.47568, 161.41096, 161.46745, 161.4061, 161.49786, 161.47142, 161.59058, 161.50833, 161.52203, 161.54617, 161.53557, 161.57367, 161.53569, 161.54568, 161.55978, 161.60565, 161.61751, 161.58444, 161.6586, 161.62756, 161.68524, 161.61127, 161.67822, 161.6719, 161.70132, 161.69109, 161.75418, 161.71866, 161.724, 161.69296, 161.69424, 161.71683, 161.74167, 161.74176, 161.66241, 161.69893, 161.70308, 161.67105, 161.68384, 161.7038, 161.6625, 161.7172, 161.67365, 161.62941, 161.64908, 161.63821, 161.62436, 161.60162, 161.52771, 161.51141, 161.55164, 161.44513, 161.46457, 161.453, 161.47284, 161.45479, 161.35713, 161.33365, 161.37032, 161.34798, 161.29514, 161.41116, 161.27205, 161.26425, 161.20894, 161.18924, 161.22144, 161.15475, 161.11172, 161.16281, 161.14911, 161.12534, 161.11978, 161.0935, 161.06187, 161.04771, 161.0462, 161.09421, 161.03497, 161.00967, 161.00421, 161.01358, 161.01381, 161.03241, 161.03638, 161.0253, 160.97531, 161.0087, 160.96869, 160.98965, 161.08568, 160.99353, 161.00476, 160.97055, 160.97638, 160.98419, 161.10065, 161.11284, 161.08484, 161.05386, 161.04941, 161.1395, 161.09294, 161.18549, 161.11472, 161.1164, 161.17914, 161.18146, 161.11316, 161.19374, 161.13983, 161.2233, 161.21043, 161.22604, 161.23526, 161.27426, 161.27034, 161.26103, 161.20586, 161.28601, 161.24744, 161.26996, 161.28589, 161.25658, 161.28366, 161.2922, 161.25638, 161.31494, 161.28693, 161.28903, 161.27094, 161.23604, 161.2701, 161.29587, 161.32518, 161.30804, 161.27957, 161.28986, 161.32634, 161.32828, 161.32526, 161.36758, 161.36252, 161.33026, 161.36514, 161.39346, 161.41035, 161.39305, 161.38188, 161.402, 161.44719, 161.42401, 161.44666, 161.46362, 161.46103, 161.50206, 161.52359, 161.50003, 161.52678, 161.54239, 161.55383, 161.59103, 161.578, 161.58667, 161.61237, 161.65247, 161.64542, 161.7222, 161.62468, 161.73853, 161.67944, 161.73906, 161.68015, 161.71082, 161.70941, 161.74205, 161.69792, 161.73051, 161.73605, 161.75494, 161.77232, 161.74443, 161.75467, 161.7533, 161.71443, 161.77881, 161.68181, 161.73566, 161.71915, 161.73082, 161.69455, 161.67221, 161.70642, 161.71222, 161.6752, 161.53836, 161.63435, 161.53725, 161.58176, 161.50037, 161.52156, 161.47571, 161.42204, 161.4537, 161.41293, 161.38367, 161.40182, 161.32573, 161.32632, 161.35268, 161.27866, 161.28384, 161.29095, 161.22388, 161.23807, 161.17897, 161.18123, 161.13568, 161.16013, 161.061, 161.08089, 161.13074, 161.12073, 161.10254, 161.08563, 161.03084, 161.05518, 161.02768, 161.04443, 161.03664, 161.01259, 161.01913, 161.04617, 161.04114, 160.99725, 161.0441, 161.04482, 161.11066, 161.04993, 161.09833, 161.0893, 161.04742, 161.08128, 161.12607, 161.1406, 161.18674, 161.12843, 161.11153, 161.22803, 161.15094, 161.15802, 161.26163, 161.20636, 161.23897, 161.24184, 161.28824, 161.30841, 161.3571, 161.33868, 161.3952, 161.32788, 161.45456, 161.34674, 161.3898, 156.59717, 84.94717, 1.0611382, 0.37883696, 0.3645335, 0.36033815, 0.35711563, 0.3877568, 0.3573911, 0.3546527, 0.35243675, 0.35070765, 0.34381977, 0.34183165, 0.3361806, 0.33374625, 0.33153695, 0.32710907, 0.3128551, 0.30228713, 0.29053688, 0.34572923, 0.33457345, 0.32621342, 0.33761114, 0.33490503, 0.32899487, 0.32308543, 0.3174308, 0.31569606, 0.31301272, 0.3103106, 0.31005394, 0.30858028, 0.30636105, 0.30095592, 0.30243757, 0.30318034, 0.30196592, 0.30170116, 0.30047238, 0.3031784, 0.3004642, 0.30194074, 0.3076095, 0.30612573, 0.30612168, 0.30881757, 0.31152564, 0.3125268, 0.3154775, 0.313989, 0.31473428, 0.31892174, 0.31917033, 0.32234502, 0.32233068, 0.32407278, 0.3275215, 0.32899022, 0.33073336, 0.33195525, 0.32898638, 0.329241, 0.3319425, 0.3334239, 0.33638102, 0.33711767, 0.33564043, 0.33859098, 0.3408134, 0.3435154, 0.34080976, 0.34081239, 0.34107506, 0.342287, 0.34228098, 0.34227288, 0.34646398, 0.34746718, 0.35016298, 0.35164642, 0.35163635, 0.35013413, 0.3513609, 0.3528455, 0.35703078, 0.35432893, 0.35432568, 0.35458487, 0.35755002, 0.3587702, 0.355807, 0.35485044, 0.35828787, 0.36125472, 0.3612547, 0.35928777, 0.35779622, 0.35752892, 0.35630476, 0.35900623, 0.35630476, 0.35826558, 0.36122835, 0.3641955, 0.36811435, 0.36811036, 0.36959416, 0.36984593, 0.3737595, 0.3722741, 0.37178394, 0.3747493, 0.37623417, 0.37697482, 0.37697136, 0.37548536, 0.37819475, 0.38386357, 0.37966788, 0.378917, 0.38039026, 0.38038826, 0.3818709, 0.38483146, 0.3872714, 0.38753062, 0.39170116, 0.39292997, 0.3909651, 0.3906957, 0.3894756, 0.3902195, 0.3917134, 0.39292294, 0.39218313, 0.3894898, 0.38947964, 0.3902215, 0.39415377, 0.3914391, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
