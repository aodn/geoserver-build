netcdf file-8.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (52 currently)
  variables:
    float LATITUDE(DEPTH=52);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=52);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=52);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=52);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=52);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=52);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815, 22200.202939814815}
TEMP =
  {16.8613, 16.8772, 16.8791, 16.8766, 16.8622, 16.8499, 16.8444, 16.8414, 16.84, 16.838, 16.837, 16.8367, 16.8362, 16.8346, 16.8325, 16.8317, 16.8302, 16.8303, 16.8296, 16.8296, 16.8282, 16.8266, 16.826, 16.8254, 16.8251, 16.8249, 16.8245, 16.8238, 16.8238, 16.8238, 16.8238, 16.8228, 16.8204, 16.8201, 16.82, 16.8189, 16.8187, 16.8191, 16.8189, 16.8185, 16.8188, 16.8186, 16.8184, 16.8181, 16.8173, 16.8169, 16.8162, 16.8152, 16.815, 16.8145, 16.8136, 16.8131}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0}
}
