netcdf file-9.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (41 currently)
  variables:
    float LATITUDE(DEPTH=41);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=41);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=41);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=41);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=41);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=41);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625, 22299.0665625}
TEMP =
  {20.4294, 20.4287, 20.4287, 20.4286, 20.4288, 20.4264, 20.4206, 20.4215, 20.4145, 20.4089, 20.4052, 20.4037, 20.4011, 20.3997, 20.3935, 20.3912, 20.3903, 20.386, 20.3808, 20.3743, 20.3659, 20.3496, 20.3333, 20.3237, 20.2974, 20.2547, 20.1979, 20.1312, 20.0671, 20.0145, 19.9862, 19.8995, 19.6887, 19.6069, 19.5718, 19.5288, 19.4958, 19.4841, 19.4714, 19.4426, 19.4243}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0}
}
