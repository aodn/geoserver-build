netcdf file-147.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (27 currently)
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875, 21801.071875}
TEMP =
  {24.6823, 24.7729, 24.7846, 24.8379, 24.837, 24.8369, 24.8378, 24.8406, 24.8419, 24.8389, 24.8373, 24.8366, 24.8356, 24.8354, 24.8353, 24.835, 24.8348, 24.8351, 24.8356, 24.836, 24.8361, 24.8362, 24.8359, 24.8356, 24.8348, 24.8338, 24.834}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835}
}
