netcdf file-10.nc {
  dimensions:
    DEPTH = 50;
  variables:
    float LATITUDE(DEPTH=50);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=50);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=50);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=50);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=50);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=50);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625, 22411.1090625}
TEMP =
  {20.5721, 20.5763, 20.5743, 20.5751, 20.5697, 20.5615, 20.5542, 20.5519, 20.555, 20.5472, 20.5427, 20.5437, 20.5439, 20.5454, 20.5436, 20.5416, 20.5322, 20.5221, 20.5163, 20.5149, 20.5111, 20.5063, 20.5017, 20.502, 20.497, 20.49, 20.484, 20.4728, 20.4638, 20.4501, 20.4442, 20.4374, 20.4281, 20.422, 20.4172, 20.4132, 20.4074, 20.3993, 20.3951, 20.3889, 20.3839, 20.3806, 20.3796, 20.3784, 20.3767, 20.3727, 20.3608, 20.3263, 20.2313, 20.1795}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0}
}
