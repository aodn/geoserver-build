netcdf file-54.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (44 currently)
  variables:
    float LATITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=44);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=44);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008, -32.000008}
LONGITUDE =
  {115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664}
TIME =
  {22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111, 22998.18298611111}
TEMP =
  {20.9662, 20.9586, 20.9508, 20.9391, 20.9341, 20.9193, 20.9019, 20.8846, 20.8591, 20.827, 20.8129, 20.7932, 20.7618, 20.7417, 20.722, 20.6517, 20.5429, 20.5017, 20.4824, 20.4764, 20.4756, 20.4752, 20.4718, 20.4701, 20.4687, 20.468, 20.465, 20.4527, 20.4481, 20.4501, 20.452, 20.4536, 20.4507, 20.4501, 20.4494, 20.4475, 20.4485, 20.4521, 20.4565, 20.4616, 20.4624, 20.4639, 20.4651, 20.47}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0}
}
