netcdf file-6.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (39 currently)
  variables:
    float LATITUDE(DEPTH=39);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=39);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=39);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=39);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=39);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=39);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926, 21995.221550925926}
TEMP =
  {19.3793, 19.2898, 19.2359, 19.2033, 19.1839, 19.1719, 19.1617, 19.148, 19.1222, 19.07, 18.9809, 18.8695, 18.7501, 18.6586, 18.5963, 18.5429, 18.5168, 18.4856, 18.4579, 18.4432, 18.434, 18.4245, 18.4126, 18.4052, 18.3991, 18.3909, 18.3779, 18.3584, 18.3157, 18.2657, 18.2242, 18.1977, 18.1712, 18.1317, 18.0813, 18.0187, 17.9469, 17.8142, 17.6666}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
