netcdf file-12.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (43 currently)
  variables:
    float LATITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=43);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=43);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815, 22613.297002314815}
TEMP =
  {18.8999, 18.9003, 18.901, 18.9033, 18.9032, 18.9033, 18.906, 18.9054, 18.9049, 18.9053, 18.9047, 18.9048, 18.9045, 18.9048, 18.9056, 18.9057, 18.9035, 18.9029, 18.9024, 18.9029, 18.9048, 18.9026, 18.903, 18.9033, 18.9053, 18.9058, 18.9, 18.881, 18.8714, 18.8702, 18.8648, 18.8495, 18.8275, 18.8065, 18.8057, 18.7978, 18.792, 18.784, 18.7754, 18.7727, 18.771, 18.7695, 18.7682}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0}
}
