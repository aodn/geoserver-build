netcdf file-106.nc {
  dimensions:
    DEPTH = 13;
  variables:
    float LATITUDE(DEPTH=13);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=13);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=13);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=13);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=13);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=13);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074, 22659.18886574074}
TEMP =
  {31.5239, 31.5229, 31.5227, 31.5231, 31.5227, 31.5223, 31.5222, 31.5223, 31.5225, 31.5225, 31.5227, 31.5229, 31.5234}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {5.966, 6.96, 7.954, 8.948, 9.943, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896}
}
