netcdf file-123.nc {
  dimensions:
    DEPTH = 22;
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111, 22988.14704861111}
TEMP =
  {32.2249, 32.2256, 32.2044, 32.1429, 32.0557, 32.0014, 31.9806, 31.9698, 31.962, 31.9534, 31.9451, 31.9354, 31.9282, 31.9244, 31.9177, 31.9124, 31.9095, 31.9073, 31.9046, 31.9007, 31.8988, 31.8986}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.885, 20.879, 21.873, 22.867}
}
