netcdf file-128.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (28 currently)
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889, 22998.02045138889}
TEMP =
  {28.2293, 28.1114, 28.0638, 28.0455, 28.0372, 28.033, 28.0323, 28.0324, 28.0313, 28.0303, 28.0301, 28.0294, 28.0282, 28.028, 28.0275, 28.0271, 28.0272, 28.0271, 28.0271, 28.0273, 28.0274, 28.0275, 28.0277, 28.0278, 28.0278, 28.0295, 28.0308, 28.0331}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
