netcdf file-112.nc {
  dimensions:
    DEPTH = 21;
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742, 22987.769803240742}
TEMP =
  {31.9955, 32.0062, 32.0053, 32.0057, 32.0059, 32.0071, 32.0069, 32.0067, 32.0075, 32.0088, 32.0096, 32.0099, 32.0097, 32.0088, 32.0067, 32.0054, 32.0051, 32.0051, 32.0047, 32.004, 32.0037}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879, 21.873}
}
