netcdf file-42.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (44 currently)
  variables:
    float LATITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=44);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=44);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074, 22485.11667824074}
TEMP =
  {19.9875, 19.9878, 19.9881, 19.988, 19.9888, 19.9886, 19.9865, 19.9864, 19.9852, 19.9847, 19.9845, 19.9844, 19.9846, 19.9848, 19.9867, 19.9875, 19.9874, 19.9794, 19.8778, 19.5925, 19.194, 19.0587, 18.9594, 18.9178, 18.9251, 18.9335, 18.9654, 18.9676, 18.9566, 18.9562, 18.9355, 18.8672, 18.8381, 18.8203, 18.8146, 18.8107, 18.8086, 18.8084, 18.8074, 18.8078, 18.8082, 18.8084, 18.8084, 18.8084}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
