netcdf file-13.nc {
  dimensions:
    DEPTH = 44;
  variables:
    float LATITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=44);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=44);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518, 22704.096331018518}
TEMP =
  {20.8474, 20.8609, 20.8662, 20.8687, 20.8716, 20.8696, 20.8662, 20.8718, 20.8732, 20.8709, 20.8709, 20.8716, 20.8738, 20.876, 20.877, 20.8771, 20.8778, 20.878, 20.8778, 20.8776, 20.8778, 20.878, 20.8778, 20.8776, 20.878, 20.8791, 20.8803, 20.8808, 20.881, 20.8805, 20.8797, 20.8783, 20.8772, 20.8781, 20.8782, 20.8739, 20.8739, 20.8726, 20.8716, 20.8695, 20.8666, 20.8635, 20.86, 20.8567}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0}
}
