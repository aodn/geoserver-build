netcdf file-86.nc {
  dimensions:
    DEPTH = 22;
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076, 23178.541886574076}
TEMP =
  {27.0709, 27.1116, 27.1104, 27.1121, 27.1127, 27.113, 27.1134, 27.1116, 27.106, 27.0992, 27.0901, 27.084, 27.0796, 27.0724, 27.07, 27.0691, 27.0662, 27.0626, 27.0596, 27.0566, 27.0536, 27.0514}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866}
}
