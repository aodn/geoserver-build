netcdf file-90.nc {
  dimensions:
    DEPTH = 22;
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298, 23178.708483796298}
TEMP =
  {27.0906, 27.0741, 27.0716, 27.0733, 27.073, 27.0774, 27.082, 27.0883, 27.093, 27.095, 27.0956, 27.0956, 27.0954, 27.0951, 27.0947, 27.0941, 27.0928, 27.0921, 27.0931, 27.0934, 27.0917, 27.0909}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.902, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866}
}
