netcdf file-153.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (23 currently)
  variables:
    float LATITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=23);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=23);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963, 22055.05650462963}
TEMP =
  {24.8092, 24.8126, 24.8014, 24.7923, 24.7894, 24.7877, 24.787, 24.7872, 24.7877, 24.7874, 24.7869, 24.7872, 24.7873, 24.7874, 24.7874, 24.7876, 24.7874, 24.7877, 24.7892, 24.7901, 24.7901, 24.7897, 24.7888}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853}
}
