netcdf IMOS_ANMN-TS_20150113T230000Z_NRSROT-ADCP_FV01_NRSROT-ADCP-1409-RDI-WHS600-44_END-20150129T030000Z_id-7740.nc {
  dimensions:
    TIME = UNLIMITED;   // (729 currently)
  variables:
    double TIME(TIME=729);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=729);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=729);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=729);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=729);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=729);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=729);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=729);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=729);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=729);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=729);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=729);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=729);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical max information has been computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :instrument = "RDI WHS600";
  :references = "http://www.imos.org.au";
  :site_code = "NRSROT";
  :platform_code = "NRSROT-ADCP";
  :deployment_code = "NRSROT-ADCP-1409";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "14263";
  :history = "2015-01-29T09:02:47Z - depthPP: Depth computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).\n2015-01-29T09:02:50Z - magneticDeclinationPP: data initially referring to magnetic North has been modified so that it now refers to true North, applying a computed magnetic declination of -1.9167degrees. NOAA\'s Geomag v7.0 software + IGRF11 model have been used to compute this value at a latitude=-31.9966degrees North, longitude=115.4157degrees East, depth=44m (instrument nominal depth) and date=2014/11/24 (date in the middle of time_coverage_start and time_coverage_end).";
  :geospatial_lat_min = -31.9966; // double
  :geospatial_lat_max = -31.9966; // double
  :geospatial_lon_min = 115.4157166667; // double
  :geospatial_lon_max = 115.4157166667; // double
  :instrument_nominal_depth = 44.0f; // float
  :site_nominal_depth = 48.0f; // float
  :geospatial_vertical_min = -0.35384676f; // float
  :geospatial_vertical_max = 41.051956f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-09-19T05:00:00Z";
  :time_deployment_end = "2015-01-28T03:00:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-29T03:00:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.979166666668, 23754.0, 23754.020833333332, 23754.041666666668, 23754.0625, 23754.083333333332, 23754.104166666668, 23754.125, 23754.145833333332, 23754.166666666668, 23754.1875, 23754.208333333332, 23754.229166666668, 23754.25, 23754.270833333332, 23754.291666666668, 23754.3125, 23754.333333333332, 23754.354166666668, 23754.375, 23754.395833333332, 23754.416666666668, 23754.4375, 23754.458333333332, 23754.479166666668, 23754.5, 23754.520833333332, 23754.541666666668, 23754.5625, 23754.583333333332, 23754.604166666668, 23754.625, 23754.645833333332, 23754.666666666668, 23754.6875, 23754.708333333332, 23754.729166666668, 23754.75, 23754.770833333332, 23754.791666666668, 23754.8125, 23754.833333333332, 23754.854166666668, 23754.875, 23754.895833333332, 23754.916666666668, 23754.9375, 23754.958333333332, 23754.979166666668, 23755.0, 23755.020833333332, 23755.041666666668, 23755.0625, 23755.083333333332, 23755.104166666668, 23755.125, 23755.145833333332, 23755.166666666668, 23755.1875, 23755.208333333332, 23755.229166666668, 23755.25, 23755.270833333332, 23755.291666666668, 23755.3125, 23755.333333333332, 23755.354166666668, 23755.375, 23755.395833333332, 23755.416666666668, 23755.4375, 23755.458333333332, 23755.479166666668, 23755.5, 23755.520833333332, 23755.541666666668, 23755.5625, 23755.583333333332, 23755.604166666668, 23755.625, 23755.645833333332, 23755.666666666668, 23755.6875, 23755.708333333332, 23755.729166666668, 23755.75, 23755.770833333332, 23755.791666666668, 23755.8125, 23755.833333333332, 23755.854166666668, 23755.875, 23755.895833333332, 23755.916666666668, 23755.9375, 23755.958333333332, 23755.979166666668, 23756.0, 23756.020833333332, 23756.041666666668, 23756.0625, 23756.083333333332, 23756.104166666668, 23756.125, 23756.145833333332, 23756.166666666668, 23756.1875, 23756.208333333332, 23756.229166666668, 23756.25, 23756.270833333332, 23756.291666666668, 23756.3125, 23756.333333333332, 23756.354166666668, 23756.375, 23756.395833333332, 23756.416666666668, 23756.4375, 23756.458333333332, 23756.479166666668, 23756.5, 23756.520833333332, 23756.541666666668, 23756.5625, 23756.583333333332, 23756.604166666668, 23756.625, 23756.645833333332, 23756.666666666668, 23756.6875, 23756.708333333332, 23756.729166666668, 23756.75, 23756.770833333332, 23756.791666666668, 23756.8125, 23756.833333333332, 23756.854166666668, 23756.875, 23756.895833333332, 23756.916666666668, 23756.9375, 23756.958333333332, 23756.979166666668, 23757.0, 23757.020833333332, 23757.041666666668, 23757.0625, 23757.083333333332, 23757.104166666668, 23757.125, 23757.145833333332, 23757.166666666668, 23757.1875, 23757.208333333332, 23757.229166666668, 23757.25, 23757.270833333332, 23757.291666666668, 23757.3125, 23757.333333333332, 23757.354166666668, 23757.375, 23757.395833333332, 23757.416666666668, 23757.4375, 23757.458333333332, 23757.479166666668, 23757.5, 23757.520833333332, 23757.541666666668, 23757.5625, 23757.583333333332, 23757.604166666668, 23757.625, 23757.645833333332, 23757.666666666668, 23757.6875, 23757.708333333332, 23757.729166666668, 23757.75, 23757.770833333332, 23757.791666666668, 23757.8125, 23757.833333333332, 23757.854166666668, 23757.875, 23757.895833333332, 23757.916666666668, 23757.9375, 23757.958333333332, 23757.979166666668, 23758.0, 23758.020833333332, 23758.041666666668, 23758.0625, 23758.083333333332, 23758.104166666668, 23758.125, 23758.145833333332, 23758.166666666668, 23758.1875, 23758.208333333332, 23758.229166666668, 23758.25, 23758.270833333332, 23758.291666666668, 23758.3125, 23758.333333333332, 23758.354166666668, 23758.375, 23758.395833333332, 23758.416666666668, 23758.4375, 23758.458333333332, 23758.479166666668, 23758.5, 23758.520833333332, 23758.541666666668, 23758.5625, 23758.583333333332, 23758.604166666668, 23758.625, 23758.645833333332, 23758.666666666668, 23758.6875, 23758.708333333332, 23758.729166666668, 23758.75, 23758.770833333332, 23758.791666666668, 23758.8125, 23758.833333333332, 23758.854166666668, 23758.875, 23758.895833333332, 23758.916666666668, 23758.9375, 23758.958333333332, 23758.979166666668, 23759.0, 23759.020833333332, 23759.041666666668, 23759.0625, 23759.083333333332, 23759.104166666668, 23759.125, 23759.145833333332, 23759.166666666668, 23759.1875, 23759.208333333332, 23759.229166666668, 23759.25, 23759.270833333332, 23759.291666666668, 23759.3125, 23759.333333333332, 23759.354166666668, 23759.375, 23759.395833333332, 23759.416666666668, 23759.4375, 23759.458333333332, 23759.479166666668, 23759.5, 23759.520833333332, 23759.541666666668, 23759.5625, 23759.583333333332, 23759.604166666668, 23759.625, 23759.645833333332, 23759.666666666668, 23759.6875, 23759.708333333332, 23759.729166666668, 23759.75, 23759.770833333332, 23759.791666666668, 23759.8125, 23759.833333333332, 23759.854166666668, 23759.875, 23759.895833333332, 23759.916666666668, 23759.9375, 23759.958333333332, 23759.979166666668, 23760.0, 23760.020833333332, 23760.041666666668, 23760.0625, 23760.083333333332, 23760.104166666668, 23760.125, 23760.145833333332, 23760.166666666668, 23760.1875, 23760.208333333332, 23760.229166666668, 23760.25, 23760.270833333332, 23760.291666666668, 23760.3125, 23760.333333333332, 23760.354166666668, 23760.375, 23760.395833333332, 23760.416666666668, 23760.4375, 23760.458333333332, 23760.479166666668, 23760.5, 23760.520833333332, 23760.541666666668, 23760.5625, 23760.583333333332, 23760.604166666668, 23760.625, 23760.645833333332, 23760.666666666668, 23760.6875, 23760.708333333332, 23760.729166666668, 23760.75, 23760.770833333332, 23760.791666666668, 23760.8125, 23760.833333333332, 23760.854166666668, 23760.875, 23760.895833333332, 23760.916666666668, 23760.9375, 23760.958333333332, 23760.979166666668, 23761.0, 23761.020833333332, 23761.041666666668, 23761.0625, 23761.083333333332, 23761.104166666668, 23761.125, 23761.145833333332, 23761.166666666668, 23761.1875, 23761.208333333332, 23761.229166666668, 23761.25, 23761.270833333332, 23761.291666666668, 23761.3125, 23761.333333333332, 23761.354166666668, 23761.375, 23761.395833333332, 23761.416666666668, 23761.4375, 23761.458333333332, 23761.479166666668, 23761.5, 23761.520833333332, 23761.541666666668, 23761.5625, 23761.583333333332, 23761.604166666668, 23761.625, 23761.645833333332, 23761.666666666668, 23761.6875, 23761.708333333332, 23761.729166666668, 23761.75, 23761.770833333332, 23761.791666666668, 23761.8125, 23761.833333333332, 23761.854166666668, 23761.875, 23761.895833333332, 23761.916666666668, 23761.9375, 23761.958333333332, 23761.979166666668, 23762.0, 23762.020833333332, 23762.041666666668, 23762.0625, 23762.083333333332, 23762.104166666668, 23762.125, 23762.145833333332, 23762.166666666668, 23762.1875, 23762.208333333332, 23762.229166666668, 23762.25, 23762.270833333332, 23762.291666666668, 23762.3125, 23762.333333333332, 23762.354166666668, 23762.375, 23762.395833333332, 23762.416666666668, 23762.4375, 23762.458333333332, 23762.479166666668, 23762.5, 23762.520833333332, 23762.541666666668, 23762.5625, 23762.583333333332, 23762.604166666668, 23762.625, 23762.645833333332, 23762.666666666668, 23762.6875, 23762.708333333332, 23762.729166666668, 23762.75, 23762.770833333332, 23762.791666666668, 23762.8125, 23762.833333333332, 23762.854166666668, 23762.875, 23762.895833333332, 23762.916666666668, 23762.9375, 23762.958333333332, 23762.979166666668, 23763.0, 23763.020833333332, 23763.041666666668, 23763.0625, 23763.083333333332, 23763.104166666668, 23763.125, 23763.145833333332, 23763.166666666668, 23763.1875, 23763.208333333332, 23763.229166666668, 23763.25, 23763.270833333332, 23763.291666666668, 23763.3125, 23763.333333333332, 23763.354166666668, 23763.375, 23763.395833333332, 23763.416666666668, 23763.4375, 23763.458333333332, 23763.479166666668, 23763.5, 23763.520833333332, 23763.541666666668, 23763.5625, 23763.583333333332, 23763.604166666668, 23763.625, 23763.645833333332, 23763.666666666668, 23763.6875, 23763.708333333332, 23763.729166666668, 23763.75, 23763.770833333332, 23763.791666666668, 23763.8125, 23763.833333333332, 23763.854166666668, 23763.875, 23763.895833333332, 23763.916666666668, 23763.9375, 23763.958333333332, 23763.979166666668, 23764.0, 23764.020833333332, 23764.041666666668, 23764.0625, 23764.083333333332, 23764.104166666668, 23764.125, 23764.145833333332, 23764.166666666668, 23764.1875, 23764.208333333332, 23764.229166666668, 23764.25, 23764.270833333332, 23764.291666666668, 23764.3125, 23764.333333333332, 23764.354166666668, 23764.375, 23764.395833333332, 23764.416666666668, 23764.4375, 23764.458333333332, 23764.479166666668, 23764.5, 23764.520833333332, 23764.541666666668, 23764.5625, 23764.583333333332, 23764.604166666668, 23764.625, 23764.645833333332, 23764.666666666668, 23764.6875, 23764.708333333332, 23764.729166666668, 23764.75, 23764.770833333332, 23764.791666666668, 23764.8125, 23764.833333333332, 23764.854166666668, 23764.875, 23764.895833333332, 23764.916666666668, 23764.9375, 23764.958333333332, 23764.979166666668, 23765.0, 23765.020833333332, 23765.041666666668, 23765.0625, 23765.083333333332, 23765.104166666668, 23765.125, 23765.145833333332, 23765.166666666668, 23765.1875, 23765.208333333332, 23765.229166666668, 23765.25, 23765.270833333332, 23765.291666666668, 23765.3125, 23765.333333333332, 23765.354166666668, 23765.375, 23765.395833333332, 23765.416666666668, 23765.4375, 23765.458333333332, 23765.479166666668, 23765.5, 23765.520833333332, 23765.541666666668, 23765.5625, 23765.583333333332, 23765.604166666668, 23765.625, 23765.645833333332, 23765.666666666668, 23765.6875, 23765.708333333332, 23765.729166666668, 23765.75, 23765.770833333332, 23765.791666666668, 23765.8125, 23765.833333333332, 23765.854166666668, 23765.875, 23765.895833333332, 23765.916666666668, 23765.9375, 23765.958333333332, 23765.979166666668, 23766.0, 23766.020833333332, 23766.041666666668, 23766.0625, 23766.083333333332, 23766.104166666668, 23766.125, 23766.145833333332, 23766.166666666668, 23766.1875, 23766.208333333332, 23766.229166666668, 23766.25, 23766.270833333332, 23766.291666666668, 23766.3125, 23766.333333333332, 23766.354166666668, 23766.375, 23766.395833333332, 23766.416666666668, 23766.4375, 23766.458333333332, 23766.479166666668, 23766.5, 23766.520833333332, 23766.541666666668, 23766.5625, 23766.583333333332, 23766.604166666668, 23766.625, 23766.645833333332, 23766.666666666668, 23766.6875, 23766.708333333332, 23766.729166666668, 23766.75, 23766.770833333332, 23766.791666666668, 23766.8125, 23766.833333333332, 23766.854166666668, 23766.875, 23766.895833333332, 23766.916666666668, 23766.9375, 23766.958333333332, 23766.979166666668, 23767.0, 23767.020833333332, 23767.041666666668, 23767.0625, 23767.083333333332, 23767.104166666668, 23767.125, 23767.145833333332, 23767.166666666668, 23767.1875, 23767.208333333332, 23767.229166666668, 23767.25, 23767.270833333332, 23767.291666666668, 23767.3125, 23767.333333333332, 23767.354166666668, 23767.375, 23767.395833333332, 23767.416666666668, 23767.4375, 23767.458333333332, 23767.479166666668, 23767.5, 23767.520833333332, 23767.541666666668, 23767.5625, 23767.583333333332, 23767.604166666668, 23767.625, 23767.645833333332, 23767.666666666668, 23767.6875, 23767.708333333332, 23767.729166666668, 23767.75, 23767.770833333332, 23767.791666666668, 23767.8125, 23767.833333333332, 23767.854166666668, 23767.875, 23767.895833333332, 23767.916666666668, 23767.9375, 23767.958333333332, 23767.979166666668, 23768.0, 23768.020833333332, 23768.041666666668, 23768.0625, 23768.083333333332, 23768.104166666668, 23768.125, 23768.145833333332, 23768.166666666668, 23768.1875, 23768.208333333332, 23768.229166666668, 23768.25, 23768.270833333332, 23768.291666666668, 23768.3125, 23768.333333333332, 23768.354166666668, 23768.375, 23768.395833333332, 23768.416666666668, 23768.4375, 23768.458333333332, 23768.479166666668, 23768.5, 23768.520833333332, 23768.541666666668, 23768.5625, 23768.583333333332, 23768.604166666668, 23768.625, 23768.645833333332, 23768.666666666668, 23768.6875, 23768.708333333332, 23768.729166666668, 23768.75, 23768.770833333332, 23768.791666666668, 23768.8125, 23768.833333333332, 23768.854166666668, 23768.875, 23768.895833333332, 23768.916666666668, 23768.9375, 23768.958333333332, 23768.979166666668, 23769.0, 23769.020833333332, 23769.041666666668, 23769.0625, 23769.083333333332, 23769.104166666668, 23769.125}
LATITUDE =-31.9966
LONGITUDE =115.4157166667
NOMINAL_DEPTH =44.0
TEMP =
  {20.1, 20.11, 20.11, 20.11, 20.12, 20.13, 20.14, 20.15, 20.15, 20.16, 20.17, 20.17, 20.18, 20.18, 20.2, 20.21, 20.21, 20.2, 20.19, 20.19, 20.19, 20.2, 20.21, 20.23, 20.25, 20.26, 20.26, 20.27, 20.27, 20.27, 20.28, 20.27, 20.28, 20.27, 20.27, 20.27, 20.27, 20.26, 20.27, 20.26, 20.25, 20.25, 20.26, 20.26, 20.26, 20.26, 20.26, 20.26, 20.25, 20.27, 20.26, 20.26, 20.26, 20.27, 20.27, 20.28, 20.29, 20.29, 20.29, 20.3, 20.3, 20.3, 20.3, 20.3, 20.3, 20.3, 20.28, 20.27, 20.24, 20.19, 20.15, 20.14, 20.13, 20.13, 20.08, 19.99, 19.9, 19.79, 19.72, 19.66, 19.58, 19.51, 19.44, 19.39, 19.35, 19.32, 19.3, 19.27, 19.25, 19.22, 19.19, 19.17, 19.14, 19.12, 19.1, 19.08, 19.06, 19.04, 19.0, 18.98, 18.96, 18.94, 18.92, 18.89, 18.88, 18.87, 18.86, 18.87, 18.86, 18.85, 18.84, 18.82, 18.82, 18.83, 18.84, 18.84, 18.84, 18.83, 18.81, 18.79, 18.78, 18.78, 18.77, 18.78, 18.77, 18.76, 18.76, 18.76, 18.74, 18.73, 18.71, 18.68, 18.64, 18.61, 18.6, 18.58, 18.56, 18.55, 18.55, 18.54, 18.54, 18.54, 18.54, 18.54, 18.55, 18.54, 18.56, 18.56, 18.55, 18.54, 18.53, 18.52, 18.54, 18.54, 18.54, 18.56, 18.57, 18.57, 18.57, 18.57, 18.56, 18.53, 18.52, 18.5, 18.47, 18.46, 18.46, 18.46, 18.46, 18.46, 18.46, 18.47, 18.46, 18.45, 18.44, 18.45, 18.45, 18.45, 18.45, 18.45, 18.46, 18.46, 18.46, 18.46, 18.46, 18.45, 18.44, 18.43, 18.42, 18.41, 18.41, 18.41, 18.41, 18.4, 18.41, 18.42, 18.42, 18.44, 18.45, 18.46, 18.46, 18.48, 18.49, 18.5, 18.51, 18.54, 18.59, 18.77, 18.91, 18.97, 18.93, 18.92, 18.94, 18.96, 18.97, 18.98, 18.98, 19.0, 19.02, 19.02, 19.0, 18.96, 18.92, 18.88, 18.87, 18.87, 18.86, 18.86, 18.87, 18.88, 18.89, 18.9, 18.91, 18.93, 18.96, 18.98, 18.98, 19.0, 19.01, 19.04, 19.06, 19.09, 19.11, 19.14, 19.17, 19.19, 19.22, 19.24, 19.27, 19.29, 19.32, 19.33, 19.35, 19.36, 19.37, 19.38, 19.39, 19.39, 19.39, 19.4, 19.41, 19.42, 19.42, 19.42, 19.44, 19.46, 19.48, 19.5, 19.52, 19.51, 19.5, 19.49, 19.48, 19.48, 19.47, 19.46, 19.46, 19.46, 19.47, 19.47, 19.47, 19.48, 19.49, 19.5, 19.51, 19.52, 19.53, 19.54, 19.56, 19.57, 19.59, 19.6, 19.6, 19.59, 19.6, 19.62, 19.63, 19.63, 19.63, 19.63, 19.63, 19.64, 19.65, 19.67, 19.67, 19.68, 19.68, 19.69, 19.7, 19.7, 19.7, 19.71, 19.73, 19.74, 19.76, 19.76, 19.75, 19.76, 19.77, 19.77, 19.79, 19.79, 19.8, 19.81, 19.82, 19.83, 19.84, 19.86, 19.87, 19.88, 19.9, 19.91, 19.92, 19.92, 19.93, 19.94, 19.95, 19.96, 19.96, 19.97, 19.98, 19.98, 19.98, 19.98, 19.98, 19.98, 19.98, 19.98, 19.99, 19.99, 19.99, 20.0, 19.99, 20.0, 20.0, 19.99, 19.99, 19.99, 19.99, 19.99, 19.99, 19.99, 19.99, 19.99, 19.99, 20.0, 20.0, 19.99, 20.0, 19.99, 20.0, 20.0, 20.0, 20.02, 20.04, 20.05, 20.04, 20.04, 20.04, 20.04, 20.05, 20.06, 20.06, 20.05, 20.05, 20.04, 20.02, 20.01, 20.01, 20.01, 20.01, 20.0, 20.0, 20.01, 20.02, 20.03, 20.02, 20.02, 20.02, 20.02, 20.02, 20.03, 20.03, 20.04, 20.04, 20.03, 20.04, 20.04, 20.06, 20.06, 20.07, 20.07, 20.06, 20.07, 20.08, 20.08, 20.08, 20.08, 20.08, 20.07, 20.08, 20.09, 20.09, 20.09, 20.08, 20.08, 20.09, 20.1, 20.1, 20.1, 20.11, 20.11, 20.12, 20.13, 20.14, 20.14, 20.15, 20.16, 20.16, 20.18, 20.19, 20.21, 20.21, 20.23, 20.23, 20.24, 20.25, 20.26, 20.26, 20.26, 20.27, 20.27, 20.28, 20.28, 20.28, 20.27, 20.27, 20.28, 20.27, 20.27, 20.28, 20.28, 20.27, 20.28, 20.28, 20.28, 20.27, 20.25, 20.25, 20.25, 20.23, 20.22, 20.21, 20.19, 20.17, 20.17, 20.17, 20.17, 20.18, 20.19, 20.18, 20.18, 20.18, 20.17, 20.15, 20.15, 20.14, 20.14, 20.14, 20.13, 20.12, 20.12, 20.11, 20.1, 20.11, 20.1, 20.11, 20.11, 20.12, 20.15, 20.16, 20.2, 20.22, 20.25, 20.25, 20.25, 20.28, 20.31, 20.32, 20.33, 20.33, 20.34, 20.26, 20.28, 20.34, 20.36, 20.32, 20.32, 20.25, 20.21, 20.17, 20.13, 20.1, 20.07, 20.06, 20.03, 20.0, 19.98, 19.97, 19.97, 19.98, 20.0, 20.02, 20.03, 20.03, 20.02, 20.02, 20.02, 19.99, 19.98, 19.98, 20.02, 20.02, 20.03, 20.01, 20.0, 19.97, 19.95, 19.93, 19.93, 19.91, 19.92, 19.91, 19.9, 19.91, 19.92, 19.93, 19.92, 19.94, 19.93, 19.95, 19.97, 19.98, 20.0, 20.01, 20.04, 20.05, 20.07, 20.09, 20.1, 20.11, 20.13, 20.16, 20.19, 20.2, 20.18, 20.19, 20.18, 20.06, 19.95, 19.82, 19.73, 19.71, 19.73, 19.74, 19.77, 19.78, 19.83, 19.88, 19.95, 20.03, 20.11, 20.13, 20.15, 20.16, 20.14, 20.12, 20.08, 20.06, 19.97, 19.94, 19.87, 19.86, 19.87, 19.86, 19.86, 19.83, 19.89, 19.92, 19.97, 20.01, 20.03, 20.06, 20.11, 20.23, 20.34, 20.45, 20.53, 20.6, 20.65, 20.62, 20.53, 20.24, 20.0, 19.84, 19.71, 19.64, 19.64, 19.62, 19.69, 19.74, 19.74, 19.75, 19.77, 19.8, 19.86, 19.92, 19.98, 19.97, 20.03, 20.05, 20.06, 19.99, 19.92, 19.89, 19.87, 19.87, 19.86, 19.82, 19.8, 19.78, 19.76, 19.74, 19.71, 19.67, 19.67, 19.67, 19.69, 19.72, 19.72, 19.75, 19.77, 19.81, 19.82, 19.86, 19.85, 19.89, 19.93, 19.99, 20.04, 20.19, 20.38, 20.34, 20.35, 20.39, 20.46, 20.45, 20.46, 20.48, 20.53, 21.45, 26.14, 26.18, 28.0, 28.25, 27.69, 27.57, 27.39, 27.29, 27.21, 27.11, 26.98, 26.85, 26.72, 26.56, 26.39, 26.2, 26.02, 25.87, 25.73, 25.63, 25.51, 25.45, 25.4, 25.35, 25.27, 25.19, 25.11, 25.03, 24.95, 24.86, 24.72, 24.51, 24.31, 24.15, 23.96, 23.77, 23.67, 23.73, 23.79, 23.83, 23.86, 23.88, 23.93, 24.02, 24.13, 24.22, 24.3, 24.3}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {40.69, 40.718, 40.712, 40.753, 40.749, 40.801, 40.824, 40.853, 40.834, 40.862, 40.864, 40.919, 40.894, 40.932, 40.944, 40.962, 40.952, 40.971, 41.016, 41.023, 40.997, 41.021, 40.997, 40.985, 41.012, 40.973, 41.006, 40.931, 40.921, 40.892, 40.882, 40.828, 40.846, 40.758, 40.792, 40.751, 40.723, 40.695, 40.703, 40.653, 40.69, 40.658, 40.648, 40.666, 40.684, 40.634, 40.658, 40.704, 40.64, 40.649, 40.697, 40.647, 40.694, 40.745, 40.799, 40.786, 40.792, 40.788, 40.826, 40.844, 40.881, 40.912, 40.905, 40.897, 40.924, 40.948, 41.023, 41.018, 41.023, 40.992, 41.011, 41.012, 41.015, 40.968, 40.979, 40.96, 40.926, 40.838, 40.827, 40.777, 40.793, 40.685, 40.694, 40.635, 40.643, 40.624, 40.605, 40.579, 40.55, 40.548, 40.534, 40.559, 40.553, 40.577, 40.567, 40.59, 40.595, 40.593, 40.611, 40.657, 40.696, 40.705, 40.709, 40.734, 40.752, 40.745, 40.752, 40.785, 40.817, 40.835, 40.819, 40.848, 40.901, 40.962, 40.976, 40.963, 40.998, 41.018, 41.03, 40.992, 41.043, 41.002, 40.988, 40.946, 40.918, 40.846, 40.859, 40.806, 40.779, 40.691, 40.629, 40.601, 40.579, 40.573, 40.513, 40.481, 40.507, 40.485, 40.475, 40.467, 40.449, 40.508, 40.491, 40.535, 40.537, 40.574, 40.564, 40.584, 40.643, 40.693, 40.689, 40.726, 40.709, 40.732, 40.724, 40.787, 40.79, 40.775, 40.797, 40.831, 40.901, 40.96, 40.978, 40.98, 41.004, 41.037, 41.096, 41.101, 41.11, 41.079, 41.076, 41.022, 40.995, 40.979, 40.927, 40.861, 40.843, 40.753, 40.704, 40.667, 40.632, 40.57, 40.539, 40.53, 40.493, 40.458, 40.447, 40.432, 40.464, 40.498, 40.55, 40.532, 40.568, 40.589, 40.638, 40.661, 40.659, 40.715, 40.688, 40.747, 40.779, 40.765, 40.794, 40.783, 40.783, 40.841, 40.799, 40.822, 40.912, 40.973, 40.973, 41.05, 41.061, 41.118, 41.128, 41.182, 41.2, 41.236, 41.195, 41.226, 41.146, 41.132, 41.103, 41.008, 40.963, 40.929, 40.855, 40.802, 40.742, 40.697, 40.654, 40.602, 40.55, 40.556, 40.532, 40.536, 40.534, 40.55, 40.578, 40.574, 40.627, 40.645, 40.697, 40.748, 40.727, 40.772, 40.803, 40.796, 40.854, 40.827, 40.823, 40.828, 40.865, 40.847, 40.882, 40.917, 40.953, 40.994, 41.039, 41.063, 41.13, 41.17, 41.19, 41.215, 41.256, 41.283, 41.277, 41.282, 41.294, 41.226, 41.241, 41.207, 41.141, 41.105, 41.052, 40.943, 40.879, 40.83, 40.779, 40.701, 40.632, 40.615, 40.585, 40.558, 40.572, 40.522, 40.559, 40.59, 40.613, 40.613, 40.7, 40.689, 40.757, 40.784, 40.814, 40.814, 40.856, 40.82, 40.861, 40.833, 40.855, 40.857, 40.869, 40.881, 40.927, 40.959, 41.003, 41.046, 41.016, 41.109, 41.17, 41.17, 41.229, 41.256, 41.264, 41.292, 41.345, 41.313, 41.28, 41.246, 41.218, 41.178, 41.1, 41.053, 40.995, 40.905, 40.882, 40.779, 40.715, 40.681, 40.636, 40.61, 40.621, 40.565, 40.579, 40.574, 40.586, 40.604, 40.659, 40.665, 40.69, 40.763, 40.786, 40.759, 40.856, 40.833, 40.884, 40.859, 40.859, 40.815, 40.783, 40.862, 40.835, 40.88, 40.862, 40.941, 40.91, 40.951, 40.973, 41.178, 41.139, 41.168, 41.133, 41.201, 41.32, 41.228, 41.321, 41.266, 41.221, 41.205, 41.182, 41.072, 41.07, 40.992, 40.86, 40.854, 40.781, 40.786, 40.709, 40.672, 40.628, 40.612, 40.644, 40.662, 40.625, 40.567, 40.642, 40.634, 40.614, 40.678, 40.695, 40.79, 40.785, 40.809, 40.82, 40.805, 40.827, 40.816, 40.823, 40.795, 40.794, 40.798, 40.861, 40.823, 40.843, 40.884, 40.953, 40.992, 41.07, 41.072, 41.075, 41.043, 41.108, 41.151, 41.101, 41.153, 41.113, 41.032, 41.113, 41.088, 41.007, 40.946, 40.945, 40.927, 40.893, 40.81, 40.735, 40.693, 40.758, 40.653, 40.644, 40.614, 40.586, 40.652, 40.606, 40.598, 40.699, 40.757, 40.743, 40.772, 40.825, 40.803, 40.758, 40.864, 40.798, 40.858, 40.905, 40.825, 40.798, 40.841, 40.807, 40.905, 40.819, 40.878, 40.836, 40.849, 40.933, 40.905, 40.983, 40.953, 41.062, 41.007, 40.991, 40.997, 41.028, 40.964, 41.015, 41.041, 40.921, 40.947, 40.934, 40.863, 40.808, 40.823, 40.797, 40.695, 40.722, 40.681, 40.67, 40.665, 40.691, 40.667, 40.712, 40.684, 40.719, 40.75, 40.786, 40.737, 40.788, 40.87, 40.894, 40.837, 40.818, 40.853, 40.881, 40.839, 40.864, 40.838, 40.822, 40.838, 40.849, 40.858, 40.881, 40.838, 40.862, 40.874, 40.913, 40.909, 40.906, 40.917, 40.963, 40.919, 40.882, 40.93, 40.884, 40.842, 40.855, 40.841, 40.865, 40.83, 40.803, 40.784, 40.698, 40.674, 40.737, 40.689, 40.651, 40.693, 40.671, 40.8, 40.727, 40.747, 40.725, 40.788, 40.845, 40.811, 40.793, 40.849, 40.826, 40.899, 40.904, 40.889, 40.933, 40.871, 40.94, 40.909, 40.921, 40.873, 40.862, 40.902, 40.961, 40.931, 40.901, 40.884, 40.902, 40.894, 40.893, 40.827, 40.874, 40.774, 40.854, 40.787, 40.828, 40.824, 40.783, 40.798, 40.796, 40.745, 40.757, 40.704, 40.683, 40.665, 40.696, 40.673, 40.692, 40.673, 40.689, 40.713, 40.733, 40.791, 40.766, 40.8, 40.837, 40.851, 40.847, 40.861, 40.867, 40.9, 40.909, 40.918, 40.914, 40.917, 40.911, 40.918, 40.919, 40.939, 40.902, 40.894, 40.915, 40.917, 40.899, 40.891, 40.892, 40.874, 40.87, 40.831, 40.815, 40.793, 40.758, 40.758, 40.754, 40.711, 40.69, 40.669, 40.648, 40.671, 40.636, 40.63, 40.625, 40.625, 40.628, 40.634, 40.655, 40.646, 40.665, 40.684, 40.71, 40.749, 40.766, 40.789, 40.824, 40.804, 40.842, 40.848, 40.893, 40.859, 40.882, 40.902, 40.891, 40.936, 40.966, 40.973, 40.953, 40.991, 40.981, 40.949, 40.953, 40.935, 40.935, 40.924, 40.907, 40.899, 40.897, 40.845, 40.836, 40.807, 40.816, 40.779, 40.715, 40.677, 40.68, 40.65, 40.637, 40.641, 40.607, 40.606, 40.574, 40.579, 40.621, 40.628, 40.661, 40.684, 40.7, 40.742, 40.76, 40.758, 40.82, 40.83, 40.852, 40.886, 31.386, -0.279, -0.281, -0.287, -0.303, -0.33, -0.331, -0.346, -0.338, -0.355, -0.336, -0.334, -0.33, -0.34, -0.32, -0.329, -0.317, -0.294, -0.294, -0.292, -0.302, -0.32, -0.319, -0.325, -0.329, -0.315, -0.309, -0.319, -0.308, -0.314, -0.283, -0.313, -0.313, -0.292, -0.298, -0.297, -0.287, -0.283, -0.285, -0.273, -0.269, -0.272, -0.268, -0.274, -0.288, -0.267, -0.285, -0.288, -0.291}
PRES_REL_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {40.402702, 40.429893, 40.423077, 40.46387, 40.457043, 40.514915, 40.53181, 40.565887, 40.54548, 40.572666, 40.576088, 40.62703, 40.60669, 40.640636, 40.65425, 40.671238, 40.66448, 40.684906, 40.729065, 40.735886, 40.708664, 40.732456, 40.708664, 40.69504, 40.7257, 40.68834, 40.718887, 40.640648, 40.630447, 40.603268, 40.593075, 40.538654, 40.55909, 40.474148, 40.501247, 40.460457, 40.43326, 40.40608, 40.416325, 40.365276, 40.402702, 40.368668, 40.365376, 40.378906, 40.39589, 40.348343, 40.368668, 40.419754, 40.355133, 40.361904, 40.406036, 40.35849, 40.406086, 40.46054, 40.511486, 40.501324, 40.501247, 40.501297, 40.53524, 40.55913, 40.593075, 40.620213, 40.61689, 40.606636, 40.63729, 40.65763, 40.735886, 40.725605, 40.735886, 40.69838, 40.71882, 40.7257, 40.725662, 40.678047, 40.688248, 40.667824, 40.64072, 40.55231, 40.542126, 40.484215, 40.504677, 40.399315, 40.406086, 40.344875, 40.3551, 40.334667, 40.321163, 40.29049, 40.26331, 40.259884, 40.249733, 40.27007, 40.263264, 40.293964, 40.280308, 40.30758, 40.307487, 40.307533, 40.32106, 40.37212, 40.409515, 40.416275, 40.423107, 40.44346, 40.46388, 40.46054, 40.46388, 40.49444, 40.528484, 40.54201, 40.531902, 40.555622, 40.610027, 40.671238, 40.68828, 40.67467, 40.708656, 40.725605, 40.739212, 40.69838, 40.75285, 40.712044, 40.695007, 40.657684, 40.6305, 40.55909, 40.572697, 40.518295, 40.48764, 40.40614, 40.34496, 40.317772, 40.29049, 40.287117, 40.229362, 40.19532, 40.21908, 40.19871, 40.1885, 40.178272, 40.16129, 40.219078, 40.20898, 40.249733, 40.2497, 40.287117, 40.280354, 40.297302, 40.3551, 40.40267, 40.406174, 40.440117, 40.423107, 40.44693, 40.43669, 40.497868, 40.504715, 40.491154, 40.511517, 40.54551, 40.610027, 40.667824, 40.688248, 40.69166, 40.71546, 40.74603, 40.80726, 40.810616, 40.81739, 40.790253, 40.783398, 40.72899, 40.708702, 40.688248, 40.63726, 40.569225, 40.552235, 40.46387, 40.419754, 40.3789, 40.344906, 40.28027, 40.253117, 40.246353, 40.208942, 40.171528, 40.161327, 40.144287, 40.178326, 40.212322, 40.26331, 40.2498, 40.280304, 40.30068, 40.35172, 40.375534, 40.37557, 40.42994, 40.399284, 40.46397, 40.48764, 40.4775, 40.504677, 40.49447, 40.49447, 40.55228, 40.511486, 40.531864, 40.620213, 40.68834, 40.68834, 40.759636, 40.76636, 40.827614, 40.841278, 40.89222, 40.909206, 40.946613, 40.90582, 40.93297, 40.8548, 40.837757, 40.814037, 40.71885, 40.67467, 40.640667, 40.56931, 40.514908, 40.453686, 40.406036, 40.365276, 40.314304, 40.26331, 40.270134, 40.2498, 40.246254, 40.249733, 40.26331, 40.290493, 40.287117, 40.34153, 40.35852, 40.406036, 40.460503, 40.43664, 40.4843, 40.51835, 40.504616, 40.562428, 40.542126, 40.53527, 40.538654, 40.572613, 40.55909, 40.593075, 40.630505, 40.661007, 40.701805, 40.74946, 40.769783, 40.83781, 40.8786, 40.895565, 40.922783, 40.963577, 40.99421, 40.987423, 40.9908, 41.00442, 40.93297, 40.95001, 40.912544, 40.854885, 40.814014, 40.759605, 40.657715, 40.58965, 40.542088, 40.48764, 40.412888, 40.344906, 40.32791, 40.297295, 40.273537, 40.283688, 40.236115, 40.27007, 40.30758, 40.324482, 40.324482, 40.41636, 40.406174, 40.467262, 40.497913, 40.52852, 40.52852, 40.56584, 40.528435, 40.569225, 40.54204, 40.56931, 40.56929, 40.579464, 40.593075, 40.63726, 40.66783, 40.708572, 40.75278, 40.729065, 40.82086, 40.8786, 40.8786, 40.932922, 40.963577, 40.973797, 41.000977, 41.051956, 41.024834, 40.987377, 40.953384, 40.92273, 40.88882, 40.814095, 40.7665, 40.708702, 40.61689, 40.593075, 40.48764, 40.42994, 40.39593, 40.348297, 40.324528, 40.33472, 40.28035, 40.29049, 40.287117, 40.30073, 40.31772, 40.37557, 40.375477, 40.402702, 40.47407, 40.501324, 40.470688, 40.56584, 40.54204, 40.59302, 40.572697, 40.572697, 40.52505, 40.49447, 40.572666, 40.54201, 40.58964, 40.572666, 40.654305, 40.620262, 40.661053, 40.68834, 40.88882, 40.851463, 40.87517, 40.84466, 40.905735, 41.02817, 40.93639, 41.028164, 40.97723, 40.933052, 40.912582, 40.89222, 40.783443, 40.78349, 40.69838, 40.57269, 40.562428, 40.491062, 40.501324, 40.423107, 40.385715, 40.33806, 40.32795, 40.35853, 40.37553, 40.338104, 40.280308, 40.355106, 40.348343, 40.32792, 40.389084, 40.40608, 40.504715, 40.49444, 40.518265, 40.528435, 40.51487, 40.542126, 40.531948, 40.53527, 40.508095, 40.504677, 40.508053, 40.569225, 40.53527, 40.552235, 40.59302, 40.661007, 40.69838, 40.78349, 40.783443, 40.786873, 40.75285, 40.81744, 40.858196, 40.810616, 40.861603, 40.824238, 40.74264, 40.824238, 40.797024, 40.715427, 40.657684, 40.657692, 40.63726, 40.60326, 40.521664, 40.446903, 40.40267, 40.474148, 40.365276, 40.35853, 40.32792, 40.30073, 40.361862, 40.317696, 40.307457, 40.40947, 40.467262, 40.457127, 40.4843, 40.538708, 40.51835, 40.474148, 40.576088, 40.508053, 40.56928, 40.61689, 40.538708, 40.508053, 40.55228, 40.514816, 40.61689, 40.531902, 40.586243, 40.548904, 40.56252, 40.644062, 40.61689, 40.691624, 40.661007, 40.773243, 40.715427, 40.701847, 40.708664, 40.739273, 40.671192, 40.725662, 40.74942, 40.630447, 40.654217, 40.6406, 40.57266, 40.521725, 40.53527, 40.511517, 40.40608, 40.433273, 40.39593, 40.385754, 40.375477, 40.40614, 40.3789, 40.423077, 40.39589, 40.433327, 40.463924, 40.501324, 40.450317, 40.501297, 40.58289, 40.60669, 40.545425, 40.531902, 40.565887, 40.593075, 40.54884, 40.576088, 40.55231, 40.531864, 40.55231, 40.56252, 40.56928, 40.593075, 40.55231, 40.572666, 40.589733, 40.62712, 40.620262, 40.613422, 40.630505, 40.67467, 40.62703, 40.593075, 40.644115, 40.59302, 40.555702, 40.56931, 40.55228, 40.572613, 40.542088, 40.51835, 40.497913, 40.41294, 40.389145, 40.450317, 40.406174, 40.36533, 40.40267, 40.382286, 40.51148, 40.43664, 40.46397, 40.436687, 40.501297, 40.555664, 40.521656, 40.504677, 40.56252, 40.53524, 40.610065, 40.613453, 40.60332, 40.644062, 40.58289, 40.650852, 40.620262, 40.630447, 40.58285, 40.572666, 40.61693, 40.671238, 40.640648, 40.610027, 40.59302, 40.61693, 40.60669, 40.60326, 40.542126, 40.589733, 40.484253, 40.562428, 40.497868, 40.538654, 40.53181, 40.49447, 40.508053, 40.504616, 40.46054, 40.467262, 40.419754, 40.3959, 40.375477, 40.409515, 40.385704, 40.40613, 40.385704, 40.406174, 40.426502, 40.443462, 40.504715, 40.474033, 40.51148, 40.545425, 40.562454, 40.55909, 40.569225, 40.576027, 40.61349, 40.620262, 40.6305, 40.623646, 40.630505, 40.62368, 40.6305, 40.62703, 40.65086, 40.61693, 40.60669, 40.63053, 40.630505, 40.610065, 40.599846, 40.603268, 40.589733, 40.58289, 40.54551, 40.52505, 40.504677, 40.474148, 40.474148, 40.467297, 40.426556, 40.402702, 40.378853, 40.365376, 40.382286, 40.348297, 40.341496, 40.338104, 40.338104, 40.33806, 40.348343, 40.368713, 40.36195, 40.375477, 40.39589, 40.419655, 40.457043, 40.474033, 40.501293, 40.53181, 40.51487, 40.555702, 40.555622, 40.60326, 40.572697, 40.593075, 40.61693, 40.599846, 40.64401, 40.674618, 40.68834, 40.661007, 40.701847, 40.688194, 40.657623, 40.661007, 40.647484, 40.647484, 40.63729, 40.62029, 40.610065, 40.606636, 40.555664, 40.548904, 40.514816, 40.531948, 40.48764, 40.42994, 40.38909, 40.38906, 40.358437, 40.348297, 40.351665, 40.317688, 40.317696, 40.287117, 40.29049, 40.33472, 40.33806, 40.375534, 40.39589, 40.41636, 40.453686, 40.474117, 40.474148, 40.528435, 40.542088, 40.56245, 40.596466, 31.161848, -0.27480936, -0.28171122, -0.2885875, -0.3023162, -0.32634673, -0.3297977, -0.3435322, -0.33321035, -0.35384676, -0.3332231, -0.33323586, -0.32634673, -0.3401122, -0.31603777, -0.32635233, -0.31259954, -0.28854355, -0.28854355, -0.28855643, -0.30232185, -0.31603777, -0.31258687, -0.3263778, -0.32635233, -0.31606886, -0.30919254, -0.31258687, -0.30574155, -0.31261796, -0.2816984, -0.30916703, -0.30916703, -0.28855643, -0.29543266, -0.29198185, -0.2885875, -0.2816984, -0.28168568, -0.27138957, -0.26450053, -0.26793864, -0.26796412, -0.27484047, -0.28512383, -0.26451328, -0.28168568, -0.28512383, -0.28510553}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
