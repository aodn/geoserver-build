netcdf file-5.nc {
  dimensions:
    DEPTH = 42;
  variables:
    float LATITUDE(DEPTH=42);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=42);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=42);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=42);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=42);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=42);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147, 21899.200335648147}
TEMP =
  {19.1879, 19.1899, 19.1866, 19.1811, 19.1774, 19.1747, 19.1707, 19.1686, 19.1676, 19.167, 19.1669, 19.1656, 19.1632, 19.1585, 19.1453, 19.1285, 19.117, 19.1035, 19.0717, 19.048, 19.0276, 19.0139, 19.0046, 18.9954, 18.9834, 18.9739, 18.9648, 18.9484, 18.9335, 18.9227, 18.9142, 18.9079, 18.9049, 18.9023, 18.8947, 18.8849, 18.8739, 18.866, 18.8612, 18.8608, 18.86, 18.8538}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0}
}
