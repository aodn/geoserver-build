netcdf file-51.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (43 currently)
  variables:
    float LATITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=43);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=43);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001}
LONGITUDE =
  {115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943, 115.41943}
TIME =
  {22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815, 22916.163252314815}
TEMP =
  {18.7759, 18.7635, 18.7595, 18.7531, 18.7474, 18.746, 18.7457, 18.7494, 18.7528, 18.7557, 18.7577, 18.7593, 18.7618, 18.7632, 18.7631, 18.7625, 18.7619, 18.7608, 18.7602, 18.7586, 18.7583, 18.7584, 18.7584, 18.7595, 18.7606, 18.7616, 18.762, 18.7631, 18.7641, 18.7652, 18.7736, 18.7929, 18.8168, 18.8269, 18.8188, 18.7864, 18.7021, 18.599, 18.5049, 18.4068, 18.338, 18.3, 18.2693}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0}
}
