netcdf file-57.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (45 currently)
  variables:
    float LATITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=45);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=45);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015, -32.000015}
LONGITUDE =
  {115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664}
TIME =
  {23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075, 23090.165949074075}
TEMP =
  {22.7697, 22.8563, 22.8169, 22.8064, 22.8037, 22.802, 22.794, 22.7892, 22.7883, 22.7882, 22.7901, 22.7955, 22.7977, 22.7945, 22.7906, 22.7903, 22.7903, 22.7922, 22.7959, 22.7918, 22.7767, 22.7689, 22.7669, 22.7664, 22.7661, 22.7637, 22.7597, 22.7584, 22.7513, 22.7449, 22.7432, 22.7402, 22.7329, 22.7356, 22.7346, 22.7349, 22.7318, 22.7266, 22.7233, 22.7161, 22.7147, 22.715, 22.7152, 22.7141, 22.714}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
