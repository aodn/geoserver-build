netcdf file-21.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (36 currently)
  variables:
    float LATITUDE(DEPTH=36);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=36);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=36);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=36);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=36);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=36);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446, 22466.156006944446}
TEMP =
  {23.7594, 23.7593, 23.7582, 23.757, 23.7576, 23.7548, 23.7462, 23.7253, 23.7258, 23.7247, 23.7157, 23.7202, 23.7128, 23.6974, 23.6946, 23.6826, 23.6705, 23.6691, 23.6795, 23.6581, 23.6457, 23.6462, 23.6178, 23.6016, 23.5895, 23.5807, 23.5697, 23.5618, 23.5575, 23.551, 23.55, 23.5502, 23.5471, 23.5444, 23.5414, 23.5403}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0}
}
