netcdf file-89.nc {
  dimensions:
    DEPTH = 22;
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889, 23178.66982638889}
TEMP =
  {27.0427, 27.0909, 27.0875, 27.0872, 27.0886, 27.0914, 27.0913, 27.0888, 27.0904, 27.0906, 27.0904, 27.0898, 27.0897, 27.0888, 27.0883, 27.0895, 27.0908, 27.0907, 27.0908, 27.0909, 27.0906, 27.0895}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866}
}
