netcdf file-114.nc {
  dimensions:
    DEPTH = 21;
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628, 22987.833067129628}
TEMP =
  {31.9525, 31.9465, 31.9511, 31.9473, 31.9497, 31.953, 31.9559, 31.9606, 31.9613, 31.9616, 31.9616, 31.9651, 31.9652, 31.9639, 31.9643, 31.965, 31.9659, 31.9661, 31.9642, 31.9644, 31.9653}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879, 21.872}
}
