netcdf IMOS_ANMN-TS_20150113T230000Z_WATR20_FV01_WATR20-1407-Seabird-SBE39-600m-temp-only-50_END-20150122T032000Z_id-7735.nc {
  dimensions:
    TIME = 1179;
  variables:
    double TIME(TIME=1179);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=1179);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=1179);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=1179);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=1179);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=1179);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=1179);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=1179);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=1179);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=1179);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=1179);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=1179);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=1179);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been filled using the DEPTH median (mooring).";
  :instrument = "Seabird         SBE39 [600m] temp only";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "3949303-4123";
  :history = "2015-01-29T06:32:00Z - depthPP: Depth computed from the 2 nearest pressure sensors available, using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 50.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = -0.16107886f; // float
  :geospatial_vertical_max = 60.850746f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-22T03:20:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.965277777777, 23753.972222222223, 23753.979166666668, 23753.98611111111, 23753.993055555555, 23754.0, 23754.006944444445, 23754.01388888889, 23754.020833333332, 23754.027777777777, 23754.034722222223, 23754.041666666668, 23754.04861111111, 23754.055555555555, 23754.0625, 23754.069444444445, 23754.07638888889, 23754.083333333332, 23754.090277777777, 23754.097222222223, 23754.104166666668, 23754.11111111111, 23754.118055555555, 23754.125, 23754.131944444445, 23754.13888888889, 23754.145833333332, 23754.152777777777, 23754.159722222223, 23754.166666666668, 23754.17361111111, 23754.180555555555, 23754.1875, 23754.194444444445, 23754.20138888889, 23754.208333333332, 23754.215277777777, 23754.222222222223, 23754.229166666668, 23754.23611111111, 23754.243055555555, 23754.25, 23754.256944444445, 23754.26388888889, 23754.270833333332, 23754.277777777777, 23754.284722222223, 23754.291666666668, 23754.29861111111, 23754.305555555555, 23754.3125, 23754.319444444445, 23754.32638888889, 23754.333333333332, 23754.340277777777, 23754.347222222223, 23754.354166666668, 23754.36111111111, 23754.368055555555, 23754.375, 23754.381944444445, 23754.38888888889, 23754.395833333332, 23754.402777777777, 23754.409722222223, 23754.416666666668, 23754.42361111111, 23754.430555555555, 23754.4375, 23754.444444444445, 23754.45138888889, 23754.458333333332, 23754.465277777777, 23754.472222222223, 23754.479166666668, 23754.48611111111, 23754.493055555555, 23754.5, 23754.506944444445, 23754.51388888889, 23754.520833333332, 23754.527777777777, 23754.534722222223, 23754.541666666668, 23754.54861111111, 23754.555555555555, 23754.5625, 23754.569444444445, 23754.57638888889, 23754.583333333332, 23754.590277777777, 23754.597222222223, 23754.604166666668, 23754.61111111111, 23754.618055555555, 23754.625, 23754.631944444445, 23754.63888888889, 23754.645833333332, 23754.652777777777, 23754.659722222223, 23754.666666666668, 23754.67361111111, 23754.680555555555, 23754.6875, 23754.694444444445, 23754.70138888889, 23754.708333333332, 23754.715277777777, 23754.722222222223, 23754.729166666668, 23754.73611111111, 23754.743055555555, 23754.75, 23754.756944444445, 23754.76388888889, 23754.770833333332, 23754.777777777777, 23754.784722222223, 23754.791666666668, 23754.79861111111, 23754.805555555555, 23754.8125, 23754.819444444445, 23754.82638888889, 23754.833333333332, 23754.840277777777, 23754.847222222223, 23754.854166666668, 23754.86111111111, 23754.868055555555, 23754.875, 23754.881944444445, 23754.88888888889, 23754.895833333332, 23754.902777777777, 23754.909722222223, 23754.916666666668, 23754.92361111111, 23754.930555555555, 23754.9375, 23754.944444444445, 23754.95138888889, 23754.958333333332, 23754.965277777777, 23754.972222222223, 23754.979166666668, 23754.98611111111, 23754.993055555555, 23755.0, 23755.006944444445, 23755.01388888889, 23755.020833333332, 23755.027777777777, 23755.034722222223, 23755.041666666668, 23755.04861111111, 23755.055555555555, 23755.0625, 23755.069444444445, 23755.07638888889, 23755.083333333332, 23755.090277777777, 23755.097222222223, 23755.104166666668, 23755.11111111111, 23755.118055555555, 23755.125, 23755.131944444445, 23755.13888888889, 23755.145833333332, 23755.152777777777, 23755.159722222223, 23755.166666666668, 23755.17361111111, 23755.180555555555, 23755.1875, 23755.194444444445, 23755.20138888889, 23755.208333333332, 23755.215277777777, 23755.222222222223, 23755.229166666668, 23755.23611111111, 23755.243055555555, 23755.25, 23755.256944444445, 23755.26388888889, 23755.270833333332, 23755.277777777777, 23755.284722222223, 23755.291666666668, 23755.29861111111, 23755.305555555555, 23755.3125, 23755.319444444445, 23755.32638888889, 23755.333333333332, 23755.340277777777, 23755.347222222223, 23755.354166666668, 23755.36111111111, 23755.368055555555, 23755.375, 23755.381944444445, 23755.38888888889, 23755.395833333332, 23755.402777777777, 23755.409722222223, 23755.416666666668, 23755.42361111111, 23755.430555555555, 23755.4375, 23755.444444444445, 23755.45138888889, 23755.458333333332, 23755.465277777777, 23755.472222222223, 23755.479166666668, 23755.48611111111, 23755.493055555555, 23755.5, 23755.506944444445, 23755.51388888889, 23755.520833333332, 23755.527777777777, 23755.534722222223, 23755.541666666668, 23755.54861111111, 23755.555555555555, 23755.5625, 23755.569444444445, 23755.57638888889, 23755.583333333332, 23755.590277777777, 23755.597222222223, 23755.604166666668, 23755.61111111111, 23755.618055555555, 23755.625, 23755.631944444445, 23755.63888888889, 23755.645833333332, 23755.652777777777, 23755.659722222223, 23755.666666666668, 23755.67361111111, 23755.680555555555, 23755.6875, 23755.694444444445, 23755.70138888889, 23755.708333333332, 23755.715277777777, 23755.722222222223, 23755.729166666668, 23755.73611111111, 23755.743055555555, 23755.75, 23755.756944444445, 23755.76388888889, 23755.770833333332, 23755.777777777777, 23755.784722222223, 23755.791666666668, 23755.79861111111, 23755.805555555555, 23755.8125, 23755.819444444445, 23755.82638888889, 23755.833333333332, 23755.840277777777, 23755.847222222223, 23755.854166666668, 23755.86111111111, 23755.868055555555, 23755.875, 23755.881944444445, 23755.88888888889, 23755.895833333332, 23755.902777777777, 23755.909722222223, 23755.916666666668, 23755.92361111111, 23755.930555555555, 23755.9375, 23755.944444444445, 23755.95138888889, 23755.958333333332, 23755.965277777777, 23755.972222222223, 23755.979166666668, 23755.98611111111, 23755.993055555555, 23756.0, 23756.006944444445, 23756.01388888889, 23756.020833333332, 23756.027777777777, 23756.034722222223, 23756.041666666668, 23756.04861111111, 23756.055555555555, 23756.0625, 23756.069444444445, 23756.07638888889, 23756.083333333332, 23756.090277777777, 23756.097222222223, 23756.104166666668, 23756.11111111111, 23756.118055555555, 23756.125, 23756.131944444445, 23756.13888888889, 23756.145833333332, 23756.152777777777, 23756.159722222223, 23756.166666666668, 23756.17361111111, 23756.180555555555, 23756.1875, 23756.194444444445, 23756.20138888889, 23756.208333333332, 23756.215277777777, 23756.222222222223, 23756.229166666668, 23756.23611111111, 23756.243055555555, 23756.25, 23756.256944444445, 23756.26388888889, 23756.270833333332, 23756.277777777777, 23756.284722222223, 23756.291666666668, 23756.29861111111, 23756.305555555555, 23756.3125, 23756.319444444445, 23756.32638888889, 23756.333333333332, 23756.340277777777, 23756.347222222223, 23756.354166666668, 23756.36111111111, 23756.368055555555, 23756.375, 23756.381944444445, 23756.38888888889, 23756.395833333332, 23756.402777777777, 23756.409722222223, 23756.416666666668, 23756.42361111111, 23756.430555555555, 23756.4375, 23756.444444444445, 23756.45138888889, 23756.458333333332, 23756.465277777777, 23756.472222222223, 23756.479166666668, 23756.48611111111, 23756.493055555555, 23756.5, 23756.506944444445, 23756.51388888889, 23756.520833333332, 23756.527777777777, 23756.534722222223, 23756.541666666668, 23756.54861111111, 23756.555555555555, 23756.5625, 23756.569444444445, 23756.57638888889, 23756.583333333332, 23756.590277777777, 23756.597222222223, 23756.604166666668, 23756.61111111111, 23756.618055555555, 23756.625, 23756.631944444445, 23756.63888888889, 23756.645833333332, 23756.652777777777, 23756.659722222223, 23756.666666666668, 23756.67361111111, 23756.680555555555, 23756.6875, 23756.694444444445, 23756.70138888889, 23756.708333333332, 23756.715277777777, 23756.722222222223, 23756.729166666668, 23756.73611111111, 23756.743055555555, 23756.75, 23756.756944444445, 23756.76388888889, 23756.770833333332, 23756.777777777777, 23756.784722222223, 23756.791666666668, 23756.79861111111, 23756.805555555555, 23756.8125, 23756.819444444445, 23756.82638888889, 23756.833333333332, 23756.840277777777, 23756.847222222223, 23756.854166666668, 23756.86111111111, 23756.868055555555, 23756.875, 23756.881944444445, 23756.88888888889, 23756.895833333332, 23756.902777777777, 23756.909722222223, 23756.916666666668, 23756.92361111111, 23756.930555555555, 23756.9375, 23756.944444444445, 23756.95138888889, 23756.958333333332, 23756.965277777777, 23756.972222222223, 23756.979166666668, 23756.98611111111, 23756.993055555555, 23757.0, 23757.006944444445, 23757.01388888889, 23757.020833333332, 23757.027777777777, 23757.034722222223, 23757.041666666668, 23757.04861111111, 23757.055555555555, 23757.0625, 23757.069444444445, 23757.07638888889, 23757.083333333332, 23757.090277777777, 23757.097222222223, 23757.104166666668, 23757.11111111111, 23757.118055555555, 23757.125, 23757.131944444445, 23757.13888888889, 23757.145833333332, 23757.152777777777, 23757.159722222223, 23757.166666666668, 23757.17361111111, 23757.180555555555, 23757.1875, 23757.194444444445, 23757.20138888889, 23757.208333333332, 23757.215277777777, 23757.222222222223, 23757.229166666668, 23757.23611111111, 23757.243055555555, 23757.25, 23757.256944444445, 23757.26388888889, 23757.270833333332, 23757.277777777777, 23757.284722222223, 23757.291666666668, 23757.29861111111, 23757.305555555555, 23757.3125, 23757.319444444445, 23757.32638888889, 23757.333333333332, 23757.340277777777, 23757.347222222223, 23757.354166666668, 23757.36111111111, 23757.368055555555, 23757.375, 23757.381944444445, 23757.38888888889, 23757.395833333332, 23757.402777777777, 23757.409722222223, 23757.416666666668, 23757.42361111111, 23757.430555555555, 23757.4375, 23757.444444444445, 23757.45138888889, 23757.458333333332, 23757.465277777777, 23757.472222222223, 23757.479166666668, 23757.48611111111, 23757.493055555555, 23757.5, 23757.506944444445, 23757.51388888889, 23757.520833333332, 23757.527777777777, 23757.534722222223, 23757.541666666668, 23757.54861111111, 23757.555555555555, 23757.5625, 23757.569444444445, 23757.57638888889, 23757.583333333332, 23757.590277777777, 23757.597222222223, 23757.604166666668, 23757.61111111111, 23757.618055555555, 23757.625, 23757.631944444445, 23757.63888888889, 23757.645833333332, 23757.652777777777, 23757.659722222223, 23757.666666666668, 23757.67361111111, 23757.680555555555, 23757.6875, 23757.694444444445, 23757.70138888889, 23757.708333333332, 23757.715277777777, 23757.722222222223, 23757.729166666668, 23757.73611111111, 23757.743055555555, 23757.75, 23757.756944444445, 23757.76388888889, 23757.770833333332, 23757.777777777777, 23757.784722222223, 23757.791666666668, 23757.79861111111, 23757.805555555555, 23757.8125, 23757.819444444445, 23757.82638888889, 23757.833333333332, 23757.840277777777, 23757.847222222223, 23757.854166666668, 23757.86111111111, 23757.868055555555, 23757.875, 23757.881944444445, 23757.88888888889, 23757.895833333332, 23757.902777777777, 23757.909722222223, 23757.916666666668, 23757.92361111111, 23757.930555555555, 23757.9375, 23757.944444444445, 23757.95138888889, 23757.958333333332, 23757.965277777777, 23757.972222222223, 23757.979166666668, 23757.98611111111, 23757.993055555555, 23758.0, 23758.006944444445, 23758.01388888889, 23758.020833333332, 23758.027777777777, 23758.034722222223, 23758.041666666668, 23758.04861111111, 23758.055555555555, 23758.0625, 23758.069444444445, 23758.07638888889, 23758.083333333332, 23758.090277777777, 23758.097222222223, 23758.104166666668, 23758.11111111111, 23758.118055555555, 23758.125, 23758.131944444445, 23758.13888888889, 23758.145833333332, 23758.152777777777, 23758.159722222223, 23758.166666666668, 23758.17361111111, 23758.180555555555, 23758.1875, 23758.194444444445, 23758.20138888889, 23758.208333333332, 23758.215277777777, 23758.222222222223, 23758.229166666668, 23758.23611111111, 23758.243055555555, 23758.25, 23758.256944444445, 23758.26388888889, 23758.270833333332, 23758.277777777777, 23758.284722222223, 23758.291666666668, 23758.29861111111, 23758.305555555555, 23758.3125, 23758.319444444445, 23758.32638888889, 23758.333333333332, 23758.340277777777, 23758.347222222223, 23758.354166666668, 23758.36111111111, 23758.368055555555, 23758.375, 23758.381944444445, 23758.38888888889, 23758.395833333332, 23758.402777777777, 23758.409722222223, 23758.416666666668, 23758.42361111111, 23758.430555555555, 23758.4375, 23758.444444444445, 23758.45138888889, 23758.458333333332, 23758.465277777777, 23758.472222222223, 23758.479166666668, 23758.48611111111, 23758.493055555555, 23758.5, 23758.506944444445, 23758.51388888889, 23758.520833333332, 23758.527777777777, 23758.534722222223, 23758.541666666668, 23758.54861111111, 23758.555555555555, 23758.5625, 23758.569444444445, 23758.57638888889, 23758.583333333332, 23758.590277777777, 23758.597222222223, 23758.604166666668, 23758.61111111111, 23758.618055555555, 23758.625, 23758.631944444445, 23758.63888888889, 23758.645833333332, 23758.652777777777, 23758.659722222223, 23758.666666666668, 23758.67361111111, 23758.680555555555, 23758.6875, 23758.694444444445, 23758.70138888889, 23758.708333333332, 23758.715277777777, 23758.722222222223, 23758.729166666668, 23758.73611111111, 23758.743055555555, 23758.75, 23758.756944444445, 23758.76388888889, 23758.770833333332, 23758.777777777777, 23758.784722222223, 23758.791666666668, 23758.79861111111, 23758.805555555555, 23758.8125, 23758.819444444445, 23758.82638888889, 23758.833333333332, 23758.840277777777, 23758.847222222223, 23758.854166666668, 23758.86111111111, 23758.868055555555, 23758.875, 23758.881944444445, 23758.88888888889, 23758.895833333332, 23758.902777777777, 23758.909722222223, 23758.916666666668, 23758.92361111111, 23758.930555555555, 23758.9375, 23758.944444444445, 23758.95138888889, 23758.958333333332, 23758.965277777777, 23758.972222222223, 23758.979166666668, 23758.98611111111, 23758.993055555555, 23759.0, 23759.006944444445, 23759.01388888889, 23759.020833333332, 23759.027777777777, 23759.034722222223, 23759.041666666668, 23759.04861111111, 23759.055555555555, 23759.0625, 23759.069444444445, 23759.07638888889, 23759.083333333332, 23759.090277777777, 23759.097222222223, 23759.104166666668, 23759.11111111111, 23759.118055555555, 23759.125, 23759.131944444445, 23759.13888888889, 23759.145833333332, 23759.152777777777, 23759.159722222223, 23759.166666666668, 23759.17361111111, 23759.180555555555, 23759.1875, 23759.194444444445, 23759.20138888889, 23759.208333333332, 23759.215277777777, 23759.222222222223, 23759.229166666668, 23759.23611111111, 23759.243055555555, 23759.25, 23759.256944444445, 23759.26388888889, 23759.270833333332, 23759.277777777777, 23759.284722222223, 23759.291666666668, 23759.29861111111, 23759.305555555555, 23759.3125, 23759.319444444445, 23759.32638888889, 23759.333333333332, 23759.340277777777, 23759.347222222223, 23759.354166666668, 23759.36111111111, 23759.368055555555, 23759.375, 23759.381944444445, 23759.38888888889, 23759.395833333332, 23759.402777777777, 23759.409722222223, 23759.416666666668, 23759.42361111111, 23759.430555555555, 23759.4375, 23759.444444444445, 23759.45138888889, 23759.458333333332, 23759.465277777777, 23759.472222222223, 23759.479166666668, 23759.48611111111, 23759.493055555555, 23759.5, 23759.506944444445, 23759.51388888889, 23759.520833333332, 23759.527777777777, 23759.534722222223, 23759.541666666668, 23759.54861111111, 23759.555555555555, 23759.5625, 23759.569444444445, 23759.57638888889, 23759.583333333332, 23759.590277777777, 23759.597222222223, 23759.604166666668, 23759.61111111111, 23759.618055555555, 23759.625, 23759.631944444445, 23759.63888888889, 23759.645833333332, 23759.652777777777, 23759.659722222223, 23759.666666666668, 23759.67361111111, 23759.680555555555, 23759.6875, 23759.694444444445, 23759.70138888889, 23759.708333333332, 23759.715277777777, 23759.722222222223, 23759.729166666668, 23759.73611111111, 23759.743055555555, 23759.75, 23759.756944444445, 23759.76388888889, 23759.770833333332, 23759.777777777777, 23759.784722222223, 23759.791666666668, 23759.79861111111, 23759.805555555555, 23759.8125, 23759.819444444445, 23759.82638888889, 23759.833333333332, 23759.840277777777, 23759.847222222223, 23759.854166666668, 23759.86111111111, 23759.868055555555, 23759.875, 23759.881944444445, 23759.88888888889, 23759.895833333332, 23759.902777777777, 23759.909722222223, 23759.916666666668, 23759.92361111111, 23759.930555555555, 23759.9375, 23759.944444444445, 23759.95138888889, 23759.958333333332, 23759.965277777777, 23759.972222222223, 23759.979166666668, 23759.98611111111, 23759.993055555555, 23760.0, 23760.006944444445, 23760.01388888889, 23760.020833333332, 23760.027777777777, 23760.034722222223, 23760.041666666668, 23760.04861111111, 23760.055555555555, 23760.0625, 23760.069444444445, 23760.07638888889, 23760.083333333332, 23760.090277777777, 23760.097222222223, 23760.104166666668, 23760.11111111111, 23760.118055555555, 23760.125, 23760.131944444445, 23760.13888888889, 23760.145833333332, 23760.152777777777, 23760.159722222223, 23760.166666666668, 23760.17361111111, 23760.180555555555, 23760.1875, 23760.194444444445, 23760.20138888889, 23760.208333333332, 23760.215277777777, 23760.222222222223, 23760.229166666668, 23760.23611111111, 23760.243055555555, 23760.25, 23760.256944444445, 23760.26388888889, 23760.270833333332, 23760.277777777777, 23760.284722222223, 23760.291666666668, 23760.29861111111, 23760.305555555555, 23760.3125, 23760.319444444445, 23760.32638888889, 23760.333333333332, 23760.340277777777, 23760.347222222223, 23760.354166666668, 23760.36111111111, 23760.368055555555, 23760.375, 23760.381944444445, 23760.38888888889, 23760.395833333332, 23760.402777777777, 23760.409722222223, 23760.416666666668, 23760.42361111111, 23760.430555555555, 23760.4375, 23760.444444444445, 23760.45138888889, 23760.458333333332, 23760.465277777777, 23760.472222222223, 23760.479166666668, 23760.48611111111, 23760.493055555555, 23760.5, 23760.506944444445, 23760.51388888889, 23760.520833333332, 23760.527777777777, 23760.534722222223, 23760.541666666668, 23760.54861111111, 23760.555555555555, 23760.5625, 23760.569444444445, 23760.57638888889, 23760.583333333332, 23760.590277777777, 23760.597222222223, 23760.604166666668, 23760.61111111111, 23760.618055555555, 23760.625, 23760.631944444445, 23760.63888888889, 23760.645833333332, 23760.652777777777, 23760.659722222223, 23760.666666666668, 23760.67361111111, 23760.680555555555, 23760.6875, 23760.694444444445, 23760.70138888889, 23760.708333333332, 23760.715277777777, 23760.722222222223, 23760.729166666668, 23760.73611111111, 23760.743055555555, 23760.75, 23760.756944444445, 23760.76388888889, 23760.770833333332, 23760.777777777777, 23760.784722222223, 23760.791666666668, 23760.79861111111, 23760.805555555555, 23760.8125, 23760.819444444445, 23760.82638888889, 23760.833333333332, 23760.840277777777, 23760.847222222223, 23760.854166666668, 23760.86111111111, 23760.868055555555, 23760.875, 23760.881944444445, 23760.88888888889, 23760.895833333332, 23760.902777777777, 23760.909722222223, 23760.916666666668, 23760.92361111111, 23760.930555555555, 23760.9375, 23760.944444444445, 23760.95138888889, 23760.958333333332, 23760.965277777777, 23760.972222222223, 23760.979166666668, 23760.98611111111, 23760.993055555555, 23761.0, 23761.006944444445, 23761.01388888889, 23761.020833333332, 23761.027777777777, 23761.034722222223, 23761.041666666668, 23761.04861111111, 23761.055555555555, 23761.0625, 23761.069444444445, 23761.07638888889, 23761.083333333332, 23761.090277777777, 23761.097222222223, 23761.104166666668, 23761.11111111111, 23761.118055555555, 23761.125, 23761.131944444445, 23761.13888888889, 23761.145833333332, 23761.152777777777, 23761.159722222223, 23761.166666666668, 23761.17361111111, 23761.180555555555, 23761.1875, 23761.194444444445, 23761.20138888889, 23761.208333333332, 23761.215277777777, 23761.222222222223, 23761.229166666668, 23761.23611111111, 23761.243055555555, 23761.25, 23761.256944444445, 23761.26388888889, 23761.270833333332, 23761.277777777777, 23761.284722222223, 23761.291666666668, 23761.29861111111, 23761.305555555555, 23761.3125, 23761.319444444445, 23761.32638888889, 23761.333333333332, 23761.340277777777, 23761.347222222223, 23761.354166666668, 23761.36111111111, 23761.368055555555, 23761.375, 23761.381944444445, 23761.38888888889, 23761.395833333332, 23761.402777777777, 23761.409722222223, 23761.416666666668, 23761.42361111111, 23761.430555555555, 23761.4375, 23761.444444444445, 23761.45138888889, 23761.458333333332, 23761.465277777777, 23761.472222222223, 23761.479166666668, 23761.48611111111, 23761.493055555555, 23761.5, 23761.506944444445, 23761.51388888889, 23761.520833333332, 23761.527777777777, 23761.534722222223, 23761.541666666668, 23761.54861111111, 23761.555555555555, 23761.5625, 23761.569444444445, 23761.57638888889, 23761.583333333332, 23761.590277777777, 23761.597222222223, 23761.604166666668, 23761.61111111111, 23761.618055555555, 23761.625, 23761.631944444445, 23761.63888888889, 23761.645833333332, 23761.652777777777, 23761.659722222223, 23761.666666666668, 23761.67361111111, 23761.680555555555, 23761.6875, 23761.694444444445, 23761.70138888889, 23761.708333333332, 23761.715277777777, 23761.722222222223, 23761.729166666668, 23761.73611111111, 23761.743055555555, 23761.75, 23761.756944444445, 23761.76388888889, 23761.770833333332, 23761.777777777777, 23761.784722222223, 23761.791666666668, 23761.79861111111, 23761.805555555555, 23761.8125, 23761.819444444445, 23761.82638888889, 23761.833333333332, 23761.840277777777, 23761.847222222223, 23761.854166666668, 23761.86111111111, 23761.868055555555, 23761.875, 23761.881944444445, 23761.88888888889, 23761.895833333332, 23761.902777777777, 23761.909722222223, 23761.916666666668, 23761.92361111111, 23761.930555555555, 23761.9375, 23761.944444444445, 23761.95138888889, 23761.958333333332, 23761.965277777777, 23761.972222222223, 23761.979166666668, 23761.98611111111, 23761.993055555555, 23762.0, 23762.006944444445, 23762.01388888889, 23762.020833333332, 23762.027777777777, 23762.034722222223, 23762.041666666668, 23762.04861111111, 23762.055555555555, 23762.0625, 23762.069444444445, 23762.07638888889, 23762.083333333332, 23762.090277777777, 23762.097222222223, 23762.104166666668, 23762.11111111111, 23762.118055555555, 23762.125, 23762.131944444445, 23762.13888888889}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =50.0
TEMP =
  {19.9658, 19.9754, 19.9121, 20.0152, 20.0693, 20.0822, 20.1438, 20.1288, 20.0913, 20.0724, 20.0674, 20.055, 20.0302, 19.9424, 19.937, 20.0016, 20.024, 20.0203, 20.0298, 20.0563, 20.0708, 20.0902, 20.0975, 20.0973, 20.0919, 20.1277, 20.197, 20.1616, 20.1621, 20.1554, 20.1454, 20.1331, 20.1093, 20.1031, 20.0993, 20.0823, 20.1269, 20.1889, 20.1984, 20.2089, 20.3057, 20.3378, 20.2908, 20.3036, 20.3232, 20.3078, 20.3216, 20.3352, 20.3361, 20.353, 20.3944, 20.384, 20.3747, 20.3898, 20.3786, 20.3605, 20.3635, 20.3806, 20.3911, 20.3557, 20.3552, 20.3736, 20.3834, 20.4421, 20.4437, 20.4596, 20.4816, 20.4182, 20.3684, 20.3372, 20.3421, 20.331, 20.314, 20.3145, 20.3483, 20.3526, 20.3068, 20.2652, 20.2519, 20.2742, 20.2923, 20.3248, 20.3698, 20.4142, 20.4465, 20.4702, 20.4847, 20.4937, 20.4904, 20.5136, 20.529, 20.5408, 20.5458, 20.5616, 20.5302, 20.5262, 20.5279, 20.5294, 20.5298, 20.533, 20.5133, 20.5074, 20.507, 20.4918, 20.524, 20.5182, 20.4933, 20.433, 20.4081, 20.4123, 20.402, 20.3994, 20.4329, 20.4356, 20.4212, 20.4183, 20.4231, 20.4186, 20.421, 20.4374, 20.4457, 20.45, 20.4556, 20.477, 20.4857, 20.4996, 20.5074, 20.5135, 20.5129, 20.5064, 20.5029, 20.5252, 20.5341, 20.5413, 20.5485, 20.5465, 20.5534, 20.5709, 20.5754, 20.5836, 20.5825, 20.5809, 20.5909, 20.5909, 20.5803, 20.5802, 20.5762, 20.5783, 20.5764, 20.5916, 20.6072, 20.6137, 20.6045, 20.6115, 20.6201, 20.6226, 20.623, 20.6223, 20.6238, 20.6228, 20.6275, 20.6313, 20.6393, 20.6632, 20.653, 20.6345, 20.6302, 20.588, 20.61, 20.5955, 20.5923, 20.6106, 20.6371, 20.6264, 20.5973, 20.5774, 20.5133, 20.4732, 20.588, 20.4608, 20.573, 20.6389, 20.6486, 20.6531, 20.6558, 20.6592, 20.639, 20.61, 20.3469, 20.3178, 20.5481, 20.5904, 20.3962, 20.4917, 20.5312, 20.6093, 20.6214, 20.6257, 20.6206, 20.6166, 20.6232, 20.5913, 20.4524, 20.5268, 20.6129, 20.6264, 20.6254, 20.4354, 20.3749, 20.3698, 20.613, 20.4134, 20.1339, 20.1039, 20.3868, 20.4175, 20.3698, 20.2354, 20.3374, 20.3469, 20.3737, 20.4105, 20.4221, 20.4189, 20.4064, 20.3808, 20.3706, 20.4122, 20.4488, 20.5906, 20.5436, 20.6416, 20.6912, 20.662, 20.515, 20.4612, 20.4689, 20.4491, 20.4467, 20.4346, 20.455, 20.4705, 20.4621, 20.4686, 20.4611, 20.4466, 20.4587, 20.4387, 20.4482, 20.4577, 20.4555, 20.4542, 20.4405, 20.1361, 20.2128, 20.2193, 20.2438, 19.9424, 19.7614, 19.624, 19.7233, 19.5555, 19.8739, 19.9609, 19.7874, 19.6814, 19.6444, 19.5983, 20.0949, 19.809, 19.842, 19.8367, 19.6493, 19.5489, 19.5186, 19.5508, 19.8982, 20.2176, 19.9996, 19.6642, 19.5396, 19.6477, 19.6633, 19.5751, 19.4597, 19.4641, 19.6075, 19.6324, 19.4974, 19.6799, 19.516, 19.4733, 19.4117, 19.4325, 19.434, 19.4326, 19.4321, 19.4334, 19.4503, 19.4629, 19.4587, 19.3665, 19.4424, 19.5034, 19.5081, 19.5208, 19.4822, 19.3285, 19.3815, 19.4054, 19.4254, 19.4369, 19.4457, 19.4394, 19.4292, 19.4157, 19.4026, 19.4493, 19.4588, 19.4798, 19.4707, 19.4773, 19.4805, 19.4617, 19.4684, 19.4568, 19.449, 19.4572, 19.4489, 19.4715, 19.4619, 19.4956, 19.529, 19.7766, 19.9387, 19.7515, 19.5039, 19.561, 19.6151, 19.6845, 19.5689, 19.6165, 19.8646, 19.9182, 20.0759, 20.0879, 20.0882, 20.0836, 20.094, 20.1198, 20.0418, 19.9254, 19.9952, 19.9667, 19.6781, 19.6884, 19.6558, 19.9974, 19.7701, 20.0255, 19.7349, 19.7334, 19.9758, 19.8422, 19.9922, 19.895, 19.8238, 19.9556, 20.3158, 20.2379, 20.2283, 20.175, 20.0816, 20.2936, 20.0184, 19.8567, 20.2941, 20.4163, 20.5319, 20.5166, 20.611, 20.6631, 20.6836, 20.7141, 20.655, 20.6929, 20.7129, 20.7174, 20.7517, 20.6408, 20.3347, 20.4377, 20.4379, 20.5396, 20.3753, 20.0812, 20.2806, 20.224, 20.0304, 20.066, 20.3012, 20.2413, 20.0427, 19.941, 19.8348, 19.9125, 19.9859, 19.9967, 20.021, 20.019, 19.9458, 19.8969, 19.9319, 19.9424, 19.9882, 20.0049, 20.1241, 20.023, 19.957, 19.9367, 19.8989, 19.8664, 19.7784, 19.7457, 19.7435, 19.4547, 19.456, 19.6068, 19.7755, 19.924, 19.9776, 19.8395, 19.7719, 19.8965, 19.8611, 19.8662, 19.9302, 19.7852, 19.7282, 19.7398, 19.4687, 19.1289, 18.9341, 19.0442, 19.194, 19.6834, 19.565, 19.5638, 19.1659, 19.247, 19.1715, 19.6769, 19.8785, 19.7315, 19.1405, 19.0005, 19.1434, 19.2358, 19.1641, 19.6498, 19.5162, 19.7137, 19.7587, 19.8174, 19.7274, 19.5083, 19.7698, 19.7962, 19.7979, 19.819, 19.8132, 19.7783, 19.7664, 19.7174, 19.7065, 19.7133, 19.6895, 19.6779, 19.6791, 19.6864, 19.6786, 19.6557, 19.6438, 19.6515, 19.6379, 19.6296, 19.9028, 20.0685, 19.9175, 19.9946, 19.9049, 19.7144, 19.6276, 19.698, 19.8532, 19.999, 19.9742, 20.0048, 20.0039, 19.9847, 19.9796, 19.9836, 20.0231, 20.0915, 20.1379, 20.172, 20.2333, 20.293, 20.3087, 20.3328, 20.3501, 20.3482, 20.3305, 20.3157, 20.2282, 20.2132, 20.2241, 20.2551, 20.2267, 20.2392, 20.2198, 20.2252, 20.2311, 20.2554, 20.2724, 20.2654, 20.2663, 20.2566, 20.2619, 20.261, 20.2633, 20.2563, 20.2035, 20.2411, 20.274, 20.2617, 20.2644, 20.2647, 20.269, 20.2682, 20.2354, 20.2557, 20.2661, 20.2502, 20.2531, 20.2642, 20.2777, 20.2682, 20.2432, 20.2036, 20.2098, 20.2154, 20.2137, 20.2654, 20.2764, 20.2674, 20.2313, 20.1554, 20.1656, 20.1698, 20.2297, 20.2345, 20.1707, 20.2087, 20.1658, 20.1971, 20.1775, 20.062, 20.0387, 20.0454, 20.0475, 20.0526, 20.0915, 20.079, 20.0809, 20.0886, 20.0884, 20.079, 20.0984, 20.1177, 20.118, 20.1315, 20.1242, 20.0997, 20.0785, 20.1231, 20.0918, 20.1593, 20.1728, 20.1697, 20.1359, 20.1156, 20.1879, 20.2047, 20.163, 20.166, 20.2086, 20.1879, 20.2047, 20.1713, 20.2277, 20.2985, 20.3147, 20.3289, 20.3328, 20.2862, 20.2282, 20.153, 20.1401, 20.1113, 20.193, 20.2054, 20.175, 20.2205, 20.3035, 20.192, 20.0252, 19.9452, 20.1357, 20.2574, 20.2024, 20.1454, 20.028, 19.9695, 19.8856, 19.8094, 19.7015, 19.5437, 19.4586, 19.567, 19.6331, 19.5283, 19.2212, 19.5599, 19.4789, 19.523, 19.5277, 19.5282, 19.6285, 19.8056, 19.5465, 19.5424, 19.6904, 19.7737, 19.8556, 19.7907, 19.983, 19.9231, 20.0243, 19.8468, 19.8884, 19.8891, 19.98, 19.7425, 19.584, 19.5256, 19.4889, 19.5028, 19.7108, 19.6279, 19.6358, 19.7478, 19.7324, 19.7023, 19.6949, 19.8125, 19.9966, 20.0743, 20.1238, 19.9872, 19.9689, 19.9505, 19.9465, 19.8714, 19.8189, 19.7947, 19.8008, 19.8055, 19.8374, 19.8492, 19.8037, 19.8187, 19.8149, 19.8449, 19.8513, 19.9043, 19.9543, 19.9054, 19.6946, 19.7908, 19.8834, 19.9688, 19.9631, 20.0316, 20.0705, 19.9713, 19.895, 19.7212, 19.7897, 19.7882, 19.7381, 19.7278, 19.7659, 19.7349, 19.7139, 19.8222, 19.9724, 20.0573, 20.1095, 20.1421, 20.1677, 20.15, 20.1244, 20.1255, 20.1113, 20.0433, 19.8414, 20.0379, 20.1856, 20.3601, 20.394, 20.3393, 20.3198, 20.315, 20.3165, 20.3024, 20.2413, 20.0903, 19.7639, 19.9563, 20.0085, 20.015, 19.9608, 19.9427, 19.8095, 19.7493, 19.7387, 19.6845, 19.7279, 19.9067, 19.7984, 19.8342, 19.8979, 19.8545, 19.7757, 19.8143, 19.7605, 19.8578, 19.9302, 19.9872, 19.9319, 20.0617, 19.9878, 19.7936, 19.8766, 19.9568, 19.9924, 19.9798, 19.8851, 19.8093, 19.7529, 19.4419, 19.207, 19.3076, 19.1062, 19.3516, 19.4542, 19.3983, 19.5957, 19.5375, 19.6826, 19.6176, 19.6178, 19.8217, 19.673, 19.6201, 19.6399, 19.6248, 19.6444, 19.7269, 19.7609, 19.7484, 19.785, 19.6958, 19.7904, 19.8792, 19.8552, 20.0611, 20.0656, 20.0125, 19.9477, 20.0665, 20.0341, 19.7682, 19.6475, 19.8132, 19.5813, 19.9293, 20.0417, 20.0045, 19.5976, 19.3984, 19.4386, 19.6506, 19.8482, 20.0873, 19.9734, 20.3735, 19.783, 19.7552, 19.5439, 19.6057, 19.8378, 19.9312, 20.0235, 20.0074, 20.1259, 20.0813, 19.9239, 19.8499, 19.8055, 19.7682, 19.7321, 19.7272, 19.5418, 19.6059, 19.8247, 20.0324, 20.103, 19.9736, 19.9351, 20.0466, 20.0406, 19.8691, 20.1088, 19.7844, 19.9889, 19.582, 19.6227, 19.6767, 19.619, 19.5574, 19.3341, 19.2985, 19.4759, 19.5157, 19.6019, 19.4448, 19.6192, 19.3836, 19.6133, 19.63, 19.4603, 19.4704, 19.4965, 19.4531, 19.4792, 19.5111, 19.6165, 19.6103, 19.57, 19.5948, 19.5721, 19.5746, 19.6097, 19.6754, 19.6288, 19.5866, 19.6572, 19.6613, 19.6968, 19.6907, 19.689, 19.655, 19.6517, 19.6523, 19.5859, 19.6406, 19.6267, 19.5902, 19.6973, 19.6068, 19.7072, 19.7773, 19.6707, 19.7331, 19.7434, 21.4347, 23.2949, 22.6727, 22.5815, 22.257, 22.3045, 22.4372, 22.052, 21.6924, 22.3532, 23.2733, 22.9586, 22.8433, 22.7781, 22.8467, 23.5441, 25.1066, 26.2321, 27.1876, 29.7536, 28.5801, 28.0474, 27.9805, 27.8337, 27.807, 27.7642, 27.7232, 27.6826, 27.636, 27.573, 27.5, 27.4241, 27.3328, 27.2371, 27.1445, 27.0553, 26.9767, 26.8952, 26.8237, 26.7485, 26.6676, 26.58, 26.4965, 26.4242, 26.3469, 26.2842, 26.2171, 26.1423, 26.065, 25.9898, 25.9179, 25.8385, 25.7595, 25.6734, 25.5891, 25.5031, 25.4188, 25.3412, 25.2573, 25.1808, 25.1075, 25.0367, 24.9633, 24.8939, 24.8275, 24.7606, 24.6974, 24.6391, 24.5803, 24.5224, 24.4682, 24.4128, 24.3588, 24.3041, 24.2486, 24.1921, 24.1308, 24.0665, 23.9957, 23.9249, 23.8509, 23.7717, 23.6913, 23.6158, 23.5491, 23.4938, 23.4446, 23.4022, 23.3648, 23.3297, 23.2945, 23.2545, 23.2069, 23.1527, 23.0958, 23.038, 22.9806, 22.9225, 22.8639, 22.8049, 22.7466, 22.6846, 22.6245, 22.5633, 22.5027, 22.4453, 22.3885, 22.3343, 22.2795, 22.2241, 22.1681, 22.1125, 22.0559, 21.9997, 21.9424, 21.8881, 21.8326, 21.7828, 21.7354, 21.6923, 21.6515, 21.6146, 21.5778, 21.545, 21.5139, 21.485, 21.4594, 21.4392, 21.4222, 21.4044, 21.3833, 21.3694, 21.3585, 21.3532, 21.3564, 21.3591, 21.3547, 21.3454, 21.3403, 21.3409, 21.3481, 21.3581, 21.3637, 21.3716, 21.3806, 21.3903, 21.4073, 21.4182, 21.44, 21.4547, 21.4591, 21.5611, 23.1601, 22.4127, 22.119, 21.9106, 22.137, 22.3236, 22.6318, 23.054, 24.9218, 25.2924, 25.2692, 25.3615, 25.5573, 25.8709, 26.0523, 26.0258, 25.9089, 25.8144, 25.7276, 25.6621, 25.6022, 25.5542, 25.539, 25.5317, 25.5113, 25.4823, 25.4546, 25.4194, 25.3876, 25.343, 25.3053, 25.3028, 25.3077, 25.3101, 25.3087, 25.309, 25.3069, 25.3048, 25.299, 25.2925, 25.2895, 25.286, 25.2832, 25.2789, 25.271, 25.2632, 25.2519, 25.2405, 25.2289, 25.2165, 25.2029, 25.1906, 25.1763, 25.1647, 25.1524, 25.1418, 25.1316, 25.1195, 25.1089, 25.099, 25.0894, 25.0804, 25.0711, 25.0626, 25.0544, 25.048, 25.0409, 25.0336, 25.0245, 25.016, 25.0073, 24.9967, 24.9856, 24.9754, 24.9653, 24.9531, 24.9427, 24.9291, 24.9171, 24.9046, 24.8922, 24.8802, 24.8691, 24.8584, 24.8493, 24.8397, 24.8306, 24.8238, 24.8154, 24.8064, 24.7968, 24.7869, 24.7775, 24.7695, 24.7625, 24.7554, 24.7487, 24.7404, 24.7328, 24.7248, 24.7159, 24.7077, 24.7024, 24.6558, 24.6104, 24.5666, 24.5169, 24.4612, 24.4057, 24.3551, 24.3119, 24.2718, 24.2329, 24.1942, 24.1555, 24.1237, 24.0994, 24.0905, 24.0955, 24.0951, 24.087, 24.0865, 24.0972, 24.1147, 24.1328, 24.1679, 24.1975, 24.221, 24.2311, 24.2541, 24.2979, 24.3253, 24.3629, 24.3959, 24.4306, 24.465, 24.4882, 24.6346, 24.7113, 24.7865}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_REL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
DEPTH =
  {60.435646, 60.13205, 60.273407, 60.16655, 60.26603, 60.378242, 60.201298, 60.321472, 60.210987, 60.141342, 60.31768, 60.139656, 60.1329, 60.207535, 60.26699, 60.243523, 60.225388, 60.265717, 60.47084, 60.34575, 60.292877, 60.403366, 60.36371, 60.39161, 60.39294, 60.368576, 60.294044, 60.295532, 60.433167, 60.29271, 60.226982, 60.190094, 60.45066, 60.54149, 60.354218, 60.439167, 60.458702, 60.54151, 60.47396, 60.444817, 60.376816, 60.422234, 60.444046, 60.3143, 60.51348, 60.4122, 60.409843, 60.45072, 60.520844, 60.510933, 60.46514, 60.430573, 60.58771, 60.681137, 60.502308, 60.52767, 60.38382, 60.381664, 60.5595, 60.4347, 60.411514, 60.440735, 60.598007, 60.47889, 60.389503, 60.501846, 60.524086, 60.529747, 60.467205, 60.45681, 60.528103, 60.584785, 60.554527, 60.603676, 60.597828, 60.469, 60.475273, 60.458878, 60.590206, 60.390125, 60.492775, 60.407784, 60.427277, 60.554005, 60.39984, 60.50753, 60.341915, 60.418495, 60.52118, 60.400436, 60.396515, 60.387886, 60.540154, 60.4254, 60.476906, 60.3916, 60.296158, 60.326702, 60.300697, 60.38947, 60.312626, 60.204338, 60.276245, 60.22467, 60.329704, 60.460632, 60.183533, 60.302094, 60.178905, 60.31668, 60.25278, 60.35476, 60.33639, 60.37001, 60.21677, 60.40721, 60.27582, 60.215755, 60.096462, 60.143333, 60.09368, 60.09375, 60.18692, 60.171265, 60.08879, 60.109432, 60.06031, 60.139427, 60.185787, 60.027863, 60.275227, 60.011353, 60.138313, 60.141846, 60.09568, 60.08461, 60.05065, 60.061935, 60.021812, 60.011696, 59.98162, 60.104683, 59.96264, 60.154995, 60.083714, 60.01133, 60.014984, 60.122158, 60.02565, 60.25369, 60.23774, 60.03012, 60.15426, 60.2067, 60.176357, 60.04984, 60.095947, 60.14096, 60.21347, 60.171627, 60.208134, 60.18627, 60.256725, 60.17572, 60.305588, 60.108246, 60.204353, 60.264, 60.389553, 60.20198, 60.223362, 60.217445, 60.192, 60.263992, 60.207123, 60.30229, 60.291267, 60.24653, 60.13347, 60.298668, 60.379772, 60.36879, 60.303856, 60.372295, 60.343136, 60.364273, 60.46663, 60.44516, 60.310364, 60.34526, 60.14746, 60.42164, 60.49775, 60.417934, 60.34993, 60.427967, 60.36561, 60.39859, 60.455933, 60.457634, 60.49372, 60.31996, 60.287575, 60.5373, 60.488132, 60.441063, 60.375004, 60.48704, 60.473007, 60.50535, 60.466724, 60.40698, 60.344193, 60.54873, 60.504753, 60.577484, 60.31276, 60.56395, 60.332535, 60.541733, 60.456287, 60.369156, 60.296715, 60.421547, 60.358578, 60.323242, 60.21151, 60.36036, 60.3695, 60.309395, 60.388123, 60.272404, 60.492577, 60.20266, 60.303646, 60.358627, 60.383926, 60.339226, 60.21762, 60.292664, 60.348824, 60.15778, 60.034676, 60.45833, 60.198906, 60.142715, 60.125084, 60.171448, 60.150238, 60.209923, 60.256645, 60.1212, 60.04589, 60.161655, 60.193665, 60.0886, 59.923454, 60.039604, 60.166885, 60.170204, 60.143753, 60.11403, 60.033493, 59.926098, 59.96354, 59.96525, 60.109825, 59.96058, 59.9879, 60.07013, 59.949104, 60.163094, 59.93563, 60.165916, 59.990097, 60.18779, 59.953377, 60.256073, 59.930183, 59.949776, 60.119274, 60.141632, 60.005066, 60.03607, 60.064842, 59.993477, 59.952778, 60.072983, 60.062813, 60.158173, 59.94042, 59.95289, 60.21029, 60.15755, 60.13939, 60.105873, 60.236107, 60.014137, 60.2154, 60.209373, 60.104942, 60.11992, 60.175655, 60.23153, 60.282738, 60.245663, 60.200146, 60.256924, 60.24115, 60.294357, 60.157715, 60.174038, 60.13703, 60.016724, 60.164684, 60.294304, 60.33403, 60.289837, 60.252914, 60.392815, 60.248817, 60.257126, 60.37681, 60.214577, 60.308628, 60.373764, 60.35775, 60.299496, 60.38698, 60.300125, 60.3229, 60.373024, 60.395805, 60.51317, 60.611153, 60.354973, 60.427956, 60.413303, 60.494923, 60.509525, 60.483185, 60.522335, 60.619736, 60.589035, 60.517555, 60.53251, 60.60115, 60.565723, 60.544067, 60.621883, 60.510193, 60.562805, 60.488907, 60.595932, 60.49578, 60.589714, 60.598354, 60.60613, 60.436646, 60.577255, 60.498432, 60.55521, 60.490833, 60.635574, 60.644188, 60.59644, 60.529133, 60.470425, 60.589294, 60.48161, 60.52629, 60.709103, 60.417793, 60.559948, 60.683754, 60.39364, 60.53219, 60.45209, 60.4223, 60.38269, 60.448746, 60.498684, 60.268333, 60.333935, 60.33587, 60.350075, 60.274784, 60.292267, 60.383545, 60.16809, 60.23844, 60.213448, 60.280754, 60.279655, 60.182423, 60.30209, 60.118713, 60.06254, 60.243126, 60.150295, 60.09621, 60.238285, 60.177208, 60.07014, 60.046135, 59.984505, 59.874756, 60.09004, 60.03858, 60.106293, 59.873684, 59.997692, 59.85024, 60.039772, 59.99733, 60.01864, 60.093243, 60.075638, 59.960537, 60.07641, 59.982605, 59.954308, 60.04532, 60.08573, 60.004036, 59.85446, 60.002968, 59.81994, 60.069748, 60.02696, 59.84942, 59.833344, 59.986702, 60.020855, 59.95242, 60.03238, 59.977047, 60.093727, 60.057686, 60.01989, 60.154327, 60.098244, 60.19219, 60.204353, 60.050415, 60.160652, 60.10813, 60.108154, 60.16492, 60.31366, 60.30345, 60.236683, 60.256096, 60.171497, 60.31196, 60.199135, 60.14756, 60.14881, 60.27697, 60.208622, 60.01654, 60.403572, 60.23073, 60.237324, 60.24127, 60.22898, 60.245277, 60.41052, 60.26648, 60.36452, 60.40783, 60.262703, 60.35198, 60.325603, 60.56411, 60.512913, 60.398476, 60.51961, 60.526817, 60.512978, 60.585365, 60.307, 60.48487, 60.507034, 60.493755, 60.453323, 60.61667, 60.667587, 60.611725, 60.715202, 60.425682, 60.58651, 60.647663, 60.581512, 60.637665, 60.541443, 60.470932, 60.78245, 60.658173, 60.713173, 60.52453, 60.817764, 60.81606, 60.56462, 60.721413, 60.742302, 60.70671, 60.745674, 60.771782, 60.549446, 60.640305, 60.62127, 60.47753, 60.69639, 60.69819, 60.632828, 60.70769, 60.66889, 60.74048, 60.569397, 60.615845, 60.69931, 60.518684, 60.524067, 60.415962, 60.42282, 60.315998, 60.55599, 60.32466, 60.40393, 60.44033, 60.320133, 60.21291, 60.217278, 60.161747, 60.237602, 60.40061, 60.177845, 60.095245, 60.26915, 60.177036, 60.208183, 60.11801, 60.16291, 59.928482, 60.103565, 60.015617, 59.994255, 59.865837, 59.938293, 60.08947, 59.847847, 59.965508, 60.174065, 59.785645, 59.874496, 60.003452, 60.022453, 60.10932, 60.065315, 59.86574, 60.03553, 59.943577, 59.9998, 60.184906, 59.784622, 60.086807, 60.034286, 60.03441, 60.078445, 60.20666, 59.953205, 60.01564, 59.968876, 60.03024, 60.02014, 60.07457, 60.259224, 60.02549, 60.06836, 60.19339, 60.018883, 60.180515, 59.97547, 60.1112, 60.07389, 60.17569, 60.144936, 60.239872, 60.35868, 60.476273, 60.26053, 60.26505, 60.310402, 60.28549, 60.191147, 60.49148, 60.234814, 60.31964, 60.44008, 60.157845, 60.232933, 60.200634, 60.494884, 60.244667, 60.20131, 60.128517, 60.42018, 60.344933, 60.382217, 60.295963, 60.19101, 60.33055, 60.360416, 60.63561, 60.550148, 60.608932, 60.537704, 60.55281, 60.577118, 60.55053, 60.622704, 60.546417, 60.312782, 60.456173, 60.380863, 60.538605, 60.511993, 60.55075, 60.465576, 60.59945, 60.546257, 60.34388, 60.56941, 60.2789, 60.51849, 60.40103, 60.55565, 60.502747, 60.558086, 60.59068, 60.543285, 60.533302, 60.470108, 60.628624, 60.68268, 60.688183, 60.581963, 60.767933, 60.577156, 60.787292, 60.713028, 60.710823, 60.64081, 60.547268, 60.606316, 60.465027, 60.63189, 60.69046, 60.54737, 60.63508, 60.5578, 60.56196, 60.80146, 60.65718, 60.604065, 60.575325, 60.573605, 60.52072, 60.572464, 60.529404, 60.27101, 60.42199, 60.283394, 60.315414, 60.39939, 60.511497, 60.40722, 60.270885, 60.13129, 60.274673, 60.33744, 60.23578, 60.450817, 60.18715, 60.154655, 60.10981, 60.164665, 60.09343, 60.024315, 60.025154, 60.171738, 59.997444, 60.158455, 60.134193, 59.942783, 59.876175, 59.946648, 59.89061, 60.159214, 59.98913, 59.97129, 59.88552, 59.920494, 60.018013, 59.98056, 59.90473, 59.931007, 59.988804, 59.863487, 59.877663, 59.84682, 60.081367, 59.927483, 59.973175, 59.847256, 59.869072, 59.862526, 60.048252, 60.006702, 60.0502, 59.983967, 59.900467, 60.016666, 60.02367, 60.338394, 60.036415, 60.152924, 60.164223, 60.116074, 60.021553, 60.284237, 60.115456, 60.263096, 60.064316, 60.19258, 60.242107, 60.18095, 60.217422, 60.317184, 60.241165, 60.379044, 60.236298, 60.131393, 60.32599, 60.234787, 60.18917, 60.214104, 60.13993, 60.377693, 60.28393, 60.307594, 60.14533, 60.171646, 60.268158, 60.309376, 60.304787, 60.227974, 60.185814, 60.215927, 60.284473, 60.25669, 60.265137, 60.33841, 60.374626, 60.35084, 60.322475, 60.427643, 60.460426, 60.31192, 60.311417, 60.33336, 60.52322, 60.258476, 60.42, 60.482727, 60.403164, 60.40894, 60.520313, 60.48017, 60.474087, 60.515648, 60.51178, 60.518425, 60.528725, 60.570213, 60.497986, 60.71336, 60.53489, 60.736412, 60.57054, 60.7219, 60.57525, 60.712807, 60.626617, 60.650135, 60.708588, 60.667522, 60.648476, 60.722237, 60.71306, 60.670677, 60.850746, 60.707626, 60.745674, 60.675247, 60.751175, 60.798927, 60.747314, 60.76325, 60.74389, 60.788124, 60.778183, 60.69449, 60.77553, 60.78778, 60.698097, 60.533104, 60.758812, 60.54036, 60.62674, 60.490604, 60.563766, 60.44809, 60.48206, 60.555744, 60.414, 60.412003, 60.410866, 60.34724, 60.309265, 60.36407, 60.32995, 60.20043, 60.353878, 60.236042, 60.307148, 60.166367, 60.16336, 60.15889, 60.15573, 59.96292, 60.026, 60.179924, 60.128334, 60.18235, 60.10413, 60.029446, 60.0802, 60.08613, 60.053864, 60.013447, 59.935562, 59.93415, 59.994476, 60.04796, 59.963463, 60.07022, 60.03749, 60.282013, 60.07699, 60.184814, 60.179977, 60.036377, 60.11467, 60.337025, 60.229523, 60.373234, 60.23093, 60.12381, 60.442635, 60.34146, 60.2153, 60.48298, 60.294556, 60.351776, 60.307014, 60.49568, 60.52083, 60.552956, 60.606247, 60.67511, 60.45436, 60.795853, 60.567104, 60.642345, 60.592148, 2.0465295, 0.9615913, -0.09517376, -0.118676536, -0.12518385, -0.12940392, -0.07796034, -0.1255115, -0.12750502, -0.12750822, -0.12557675, -0.13245988, -0.12557994, -0.12748753, -0.13435961, -0.13131075, -0.13131075, -0.1351213, -0.13894132, -0.16107886, 0.06204779, 0.049631868, 0.044288434, -0.053108588, 0.05915091, 0.05610949, 0.05610949, 0.052685075, 0.054602608, 0.05269544, 0.050771557, 0.052689046, 0.05269225, 0.05269225, 0.048868388, 0.048865102, 0.048862018, 0.040828094, 0.042745583, 0.040828116, 0.048869133, 0.040828116, 0.040824905, 0.04886192, 0.048862018, 0.04886201, 0.05077237, 0.05268906, 0.050781876, 0.050775565, 0.05076836, 0.05077555, 0.05268906, 0.050771557, 0.05459941, 0.056112606, 0.05418879, 0.056109387, 0.056102242, 0.054188777, 0.056106288, 0.05610949, 0.054188784, 0.05609903, 0.056099135, 0.056099128, 0.056099128, 0.056109477, 0.056099143, 0.05610222, 0.05800951, 0.05610541, 0.056109484, 0.054188784, 0.05609903, 0.056102227, 0.056102227, 0.05801263, 0.056102324, 0.058012623, 0.058015812, 0.058012705, 0.05800545, 0.06297395, 0.06297715, 0.06183972, 0.06298034, 0.059929367, 0.061063673, 0.058015805, 0.05992618, 0.059929367, 0.056108605, 0.05800951, 0.058015805, 0.058015812, 0.056102324, 0.056099128, 0.058012623, 0.056102324, 0.058012623, 0.056102324, 0.058012623, 0.058012705, 0.058015805, 0.06488432, 0.06489068, 0.06489068, 0.06297, 0.06679061, 0.06679699, 0.06487629, 0.064880356, 0.0648731, 0.064873084, 0.064880356, 0.0648731, 0.066793784, 0.06870736, 0.07291339, 0.06678666, 0.06678666, 0.07290709, 0.07290708, 0.07289983, 0.07672367, 0.07481658, 0.0782305, 0.078640364, 0.07673012, 0.07864037, 0.07673012, 0.07672692, 0.07673004, 0.0801544, 0.080157585, 0.07673324, 0.07673005, 0.07824407, 0.08206477, 0.080150425, 0.0839783, 0.08015362, 0.08014722, 0.08206794, 0.08207114, 0.080150425, 0.0820576, 0.082071126, 0.08206081, 0.0020496126, -0.1293616, -0.121768996, -0.13472047, -0.14806849, -0.12712488, -0.12708987, -0.13321358, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
