netcdf file-30.nc {
  dimensions:
    DEPTH = 45;
  variables:
    float LATITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=45);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=45);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=45);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=45);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592, 22058.183217592592}
TEMP =
  {21.3311, 21.328, 21.3276, 21.3263, 21.3187, 21.3096, 21.3034, 21.3012, 21.3008, 21.3015, 21.3018, 21.3012, 21.3006, 21.3017, 21.302, 21.3017, 21.3007, 21.2998, 21.2996, 21.2994, 21.2992, 21.2993, 21.2996, 21.2994, 21.2978, 21.296, 21.2907, 21.2709, 21.2554, 21.2491, 21.2356, 21.2091, 21.1157, 21.0439, 20.9467, 20.8545, 20.6814, 20.3281, 19.9733, 19.71, 19.6167, 19.5785, 19.5435, 19.5213, 19.51}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0}
}
