netcdf file-55.nc {
  dimensions:
    DEPTH = 41;
  variables:
    float LATITUDE(DEPTH=41);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=41);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=41);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=41);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=41);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=41);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084}
LONGITUDE =
  {115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664, 115.416664}
TIME =
  {23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963, 23035.107025462963}
TEMP =
  {22.486, 22.4739, 22.4556, 22.4554, 22.4542, 22.4531, 22.4516, 22.45, 22.4493, 22.4461, 22.4369, 22.4401, 22.4459, 22.4362, 22.4284, 22.4208, 22.4115, 22.4113, 22.4122, 22.4094, 22.4071, 22.4054, 22.4018, 22.3958, 22.3873, 22.3821, 22.3741, 22.3721, 22.3574, 22.3463, 22.3415, 22.3081, 22.2638, 22.0445, 21.558, 21.2617, 21.2275, 21.1655, 20.9912, 21.0157, 20.9803}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0}
}
