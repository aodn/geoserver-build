netcdf file-148.nc {
  dimensions:
    DEPTH = 27;
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889, 21876.08638888889}
TEMP =
  {27.1812, 27.1572, 27.0985, 27.0208, 26.95, 26.8986, 26.8657, 26.8425, 26.8287, 26.8194, 26.8139, 26.8097, 26.8048, 26.7993, 26.7947, 26.7914, 26.7893, 26.7882, 26.7869, 26.7849, 26.7831, 26.7827, 26.7827, 26.7824, 26.7816, 26.7811, 26.7817}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
