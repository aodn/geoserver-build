netcdf file-28.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (50 currently)
  variables:
    float LATITUDE(DEPTH=50);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=50);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=50);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=50);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=50);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=50);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222, 23139.11565972222}
TEMP =
  {22.8816, 30.2424, 27.2831, 27.28, 27.2775, 27.2735, 27.271, 27.2713, 27.27, 27.2692, 27.2689, 27.2662, 27.2641, 27.2642, 27.2638, 27.2629, 27.2631, 27.2633, 27.263, 27.2622, 27.2656, 27.2678, 27.2739, 27.2766, 27.251, 27.2279, 27.2023, 27.1896, 27.1805, 27.1643, 27.1435, 27.1435, 27.1542, 27.1654, 27.1672, 27.1642, 27.1623, 27.1539, 27.131, 27.1167, 27.1123, 27.1088, 27.1005, 27.0792, 27.0596, 27.0392, 27.0271, 27.0129, 26.9954, 26.9866}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0}
}
