netcdf file-50.nc {
  dimensions:
    DEPTH = 46;
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185, 22853.10278935185}
TEMP =
  {20.2453, 20.2463, 20.2495, 20.2504, 20.2509, 20.2508, 20.2497, 20.2481, 20.2467, 20.2484, 20.2497, 20.2494, 20.2478, 20.246, 20.2441, 20.2439, 20.2457, 20.2467, 20.2468, 20.2482, 20.2476, 20.246, 20.2452, 20.2462, 20.2453, 20.2454, 20.2472, 20.246, 20.2425, 20.2365, 20.226, 20.212, 20.2072, 20.2044, 20.2, 20.1937, 20.1855, 20.1676, 20.1397, 20.1394, 20.1155, 20.0762, 20.0512, 20.0453, 20.0421, 99999.0}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
