netcdf file-35.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (46 currently)
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125, 22242.148125}
TEMP =
  {21.104, 21.0543, 20.9429, 20.8039, 20.7662, 20.7561, 20.7471, 20.7357, 20.7313, 20.7261, 20.7248, 20.715, 20.6956, 20.6782, 20.6734, 20.6725, 20.6707, 20.6622, 20.6559, 20.652, 20.6497, 20.6491, 20.6474, 20.6468, 20.6468, 20.6447, 20.638, 20.6275, 20.619, 20.6146, 20.6147, 20.6098, 20.6087, 20.6081, 20.6076, 20.6066, 20.6057, 20.606, 20.6061, 20.6059, 20.607, 20.6072, 20.6091, 20.6083, 20.6035, 20.6006}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
