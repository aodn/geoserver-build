netcdf file-32.nc {
  dimensions:
    DEPTH = 46;
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963, 22122.31681712963}
TEMP =
  {20.5913, 20.5934, 20.5936, 20.5923, 20.5915, 20.5907, 20.5902, 20.5895, 20.5894, 20.5887, 20.5879, 20.5868, 20.5864, 20.5834, 20.5768, 20.571, 20.5706, 20.5636, 20.5378, 20.5079, 20.488, 20.4838, 20.4828, 20.4798, 20.4767, 20.4707, 20.4616, 20.4547, 20.446, 20.4366, 20.4275, 20.4184, 20.4145, 20.4143, 20.4141, 20.4139, 20.413, 20.4108, 20.4074, 20.4034, 20.4007, 20.3933, 20.3815, 20.3629, 20.3515, 20.3412}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
