netcdf file-26.nc {
  dimensions:
    DEPTH = 51;
  variables:
    float LATITUDE(DEPTH=51);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=51);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=51);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=51);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=51);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=51);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865}
LONGITUDE =
  {113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666, 113.94666}
TIME =
  {22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446, 22956.183506944446}
TEMP =
  {23.0447, 23.0552, 23.0465, 23.0202, 22.9997, 22.9917, 22.9598, 22.9346, 22.9274, 22.9269, 22.9296, 22.9278, 22.921, 22.9173, 22.9163, 22.9176, 22.9171, 22.9157, 22.9149, 22.9142, 22.9141, 22.913, 22.911, 22.9083, 22.9091, 22.9073, 22.9055, 22.903, 22.8947, 22.8808, 22.8484, 22.8027, 22.7368, 22.6865, 22.6094, 22.5609, 22.5385, 22.5147, 22.4878, 22.4548, 22.4385, 22.4107, 22.3942, 22.3631, 22.326, 22.3131, 22.2911, 22.2617, 22.2388, 22.2211, 22.183}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0}
}
