netcdf file-87.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185, 23178.585810185185}
TEMP =
  {27.0847, 27.0942, 27.0982, 27.0983, 27.1038, 27.1079, 27.1082, 27.1075, 27.1102, 27.1102, 27.11, 27.1095, 27.1095, 27.1063, 27.1019, 27.1035, 27.1042, 27.1053, 27.1072, 27.1075, 27.1026}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872}
}
