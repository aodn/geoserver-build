netcdf file-2.nc {
  dimensions:
    DEPTH = 48;
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297, -33.93297}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816, 21681.371689814816}
TEMP =
  {19.2095, 19.2089, 19.2063, 19.2054, 19.2049, 19.2046, 19.2044, 19.2044, 19.2044, 19.2042, 19.2038, 19.2025, 19.2011, 19.2005, 19.2005, 19.2009, 19.2014, 19.2008, 19.1979, 19.1937, 19.1887, 19.1836, 19.1758, 19.1679, 19.1581, 19.1441, 19.1299, 19.116, 19.103, 19.0894, 19.08, 19.0753, 19.0696, 19.0634, 19.0598, 19.0575, 19.0561, 19.0531, 19.051, 19.0502, 19.0502, 19.0494, 19.0449, 19.0374, 19.0274, 19.0164, 19.0, 18.9474}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
