netcdf file-23.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (48 currently)
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815, 22701.07002314815}
TEMP =
  {27.0586, 27.053, 27.0539, 27.0522, 27.0505, 27.0494, 27.0505, 27.0508, 27.0507, 27.0479, 27.0436, 27.0424, 27.0429, 27.0452, 27.0442, 27.0438, 27.0423, 27.0464, 27.0473, 27.0466, 27.0245, 27.0034, 26.9964, 26.9925, 26.9853, 26.9635, 26.9411, 26.9232, 26.8951, 26.8724, 26.8704, 26.8618, 26.8328, 26.7876, 26.7688, 26.731, 26.7152, 26.6837, 26.6591, 26.647, 26.6409, 26.6258, 26.6107, 26.5904, 26.5714, 26.5565, 26.5326, 26.4759}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
