netcdf file-52.nc {
  dimensions:
    DEPTH = 46;
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084, -32.000084}
LONGITUDE =
  {115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334, 115.419334}
TIME =
  {22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482, 22937.095231481482}
TEMP =
  {19.591, 19.6131, 19.5926, 19.5926, 19.5887, 19.5811, 19.5788, 19.5736, 19.5654, 19.5545, 19.5445, 19.5386, 19.5352, 19.5337, 19.5312, 19.5261, 19.5237, 19.5213, 19.5184, 19.5159, 19.5141, 19.5119, 19.5092, 19.5067, 19.5051, 19.5043, 19.5032, 19.5014, 19.4921, 19.4599, 19.4305, 19.4093, 19.3924, 19.3813, 19.372, 19.3469, 19.3186, 19.279, 19.2111, 19.183, 19.1723, 19.1676, 19.1564, 19.1481, 19.1451, 19.1437}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
