netcdf file-74.nc {
  dimensions:
    DEPTH = 47;
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073, 22769.226886574073}
TEMP =
  {23.249874, 23.252012, 23.254436, 23.264294, 23.307648, 23.375929, 23.383356, 23.38347, 23.38232, 23.381424, 23.381363, 23.380163, 23.379105, 23.379301, 23.378382, 23.37747, 23.376995, 23.376587, 23.376596, 23.377134, 23.377392, 23.377083, 23.364462, 23.35621, 23.330223, 23.293877, 23.264809, 23.218018, 23.136198, 23.08166, 22.98042, 22.923098, 22.620842, 22.174068, 22.092695, 22.024578, 21.995972, 21.996487, 21.989521, 21.995886, 21.990261, 21.986275, 21.985533, 21.985922, 21.986, 21.985708, 21.986115}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
