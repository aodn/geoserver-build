netcdf file-20.nc {
  dimensions:
    DEPTH = 53;
  variables:
    float LATITUDE(DEPTH=53);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=53);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=53);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=53);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=53);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=53);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87, -21.87}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147, 22319.125648148147}
TEMP =
  {29.2079, 29.1446, 29.0998, 29.0657, 29.0648, 29.0654, 29.0609, 29.0587, 29.0343, 28.9512, 28.9148, 28.8626, 28.7622, 28.6915, 28.6692, 28.6632, 28.6566, 28.6573, 28.6583, 28.6531, 28.6482, 28.6488, 28.6508, 28.6513, 28.65, 28.6518, 28.6528, 28.6464, 28.64, 28.6383, 28.6383, 28.6372, 28.6369, 28.6361, 28.635, 28.6338, 28.6323, 28.6298, 28.624, 28.6145, 28.5831, 28.5654, 28.567, 28.5648, 28.5633, 28.5636, 28.5634, 28.5642, 28.5639, 28.5573, 28.5475, 28.5436, 99999.0}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0, 53.0}
}
