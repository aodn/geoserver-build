netcdf file-113.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963, 22987.81181712963}
TEMP =
  {31.9614, 31.9532, 31.9579, 31.9624, 31.9658, 31.967, 31.9674, 31.9681, 31.968, 31.9671, 31.9673, 31.9696, 31.9731, 31.9734, 31.9704, 31.9702, 31.9718, 31.9751, 31.9768, 31.9772, 31.9772}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.891, 19.884, 20.878, 21.873}
}
