netcdf file-154.nc {
  dimensions:
    DEPTH = 14;
  variables:
    float LATITUDE(DEPTH=14);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=14);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=14);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=14);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=14);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=14);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963, 22124.07400462963}
TEMP =
  {23.3512, 23.3381, 23.3261, 23.3162, 23.309, 23.3055, 23.3028, 23.3008, 23.2981, 23.2958, 23.2949, 23.2936, 23.2927, 23.2917}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853}
}
