netcdf file-40.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (48 currently)
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111, 22426.17423611111}
TEMP =
  {22.2584, 22.258, 22.2573, 22.2573, 22.2572, 22.2518, 22.2522, 22.2515, 22.2496, 22.2504, 22.2474, 22.2355, 22.1811, 22.1299, 22.0569, 21.9932, 21.9562, 21.9331, 21.8539, 21.7571, 21.7123, 21.7078, 21.7057, 21.6955, 21.6924, 21.6914, 21.6418, 21.599, 21.5829, 21.5794, 21.5764, 21.5814, 21.588, 21.5849, 21.5853, 21.5779, 21.5702, 21.5719, 21.573, 21.5674, 21.5669, 21.5696, 21.5708, 21.5744, 21.5712, 21.566, 21.5672, 21.568}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0}
}
