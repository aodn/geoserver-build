netcdf file-27.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (48 currently)
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865, -21.865}
LONGITUDE =
  {113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95, 113.95}
TIME =
  {23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852, 23050.07070601852}
TEMP =
  {28.8229, 28.7944, 28.777, 28.7546, 28.7448, 28.7406, 28.7305, 28.7366, 28.7284, 28.7123, 28.6671, 28.6508, 28.6463, 28.6429, 28.6361, 28.6271, 28.6122, 28.5925, 28.5838, 28.5704, 28.5613, 28.5571, 28.5549, 28.5514, 28.5467, 28.5447, 28.5446, 28.5449, 28.544, 28.5433, 28.5449, 28.546, 28.5455, 28.5457, 28.5447, 28.5441, 28.5432, 28.5427, 28.5429, 28.5434, 28.5438, 28.5437, 28.5438, 28.5435, 28.5448, 28.5457, 28.5432, 28.5289}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0}
}
