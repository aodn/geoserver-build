netcdf file-7.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (43 currently)
  variables:
    float LATITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=43);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=43);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625, 22094.2915625}
TEMP =
  {17.5729, 17.5779, 17.5805, 17.586, 17.5826, 17.5837, 17.5863, 17.5858, 17.585, 17.5829, 17.5816, 17.5799, 17.5811, 17.583, 17.5826, 17.5821, 17.5823, 17.5852, 17.5868, 17.5839, 17.5819, 17.5841, 17.5822, 17.5818, 17.5808, 17.5828, 17.5845, 17.5861, 17.5855, 17.5856, 17.5842, 17.5766, 17.5693, 17.5683, 17.568, 17.5652, 17.5649, 17.5655, 17.5666, 17.5694, 17.5723, 17.5704, 17.5679}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0}
}
