netcdf file-75.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (47 currently)
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001, -32.0001}
LONGITUDE =
  {115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41, 115.41}
TIME =
  {22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705, 22881.169016203705}
TEMP =
  {19.343336, 19.343801, 19.340683, 19.338066, 19.331566, 19.330286, 19.330576, 19.331078, 19.330864, 19.329344, 19.326786, 19.324423, 19.32221, 19.32055, 19.31656, 19.316135, 19.315006, 19.309643, 19.301462, 19.29926, 19.295914, 19.290369, 19.281883, 19.269358, 19.191082, 19.17605, 19.14355, 19.113615, 19.0534, 19.01598, 18.934277, 18.929686, 18.929865, 18.93071, 18.928707, 18.929838, 18.927288, 18.921858, 18.914875, 18.912733, 18.90551, 18.891312, 18.890217, 18.885511, 18.88842, 18.891449, 18.89273}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
