netcdf file-39.nc {
  dimensions:
    DEPTH = 49;
  variables:
    float LATITUDE(DEPTH=49);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=49);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=49);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=49);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=49);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=49);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928, 22362.180613425928}
TEMP =
  {24.1398, 24.1049, 24.0978, 24.0979, 23.9925, 23.8578, 23.8154, 23.8239, 23.7982, 23.7816, 23.7705, 23.7655, 23.7619, 23.7601, 23.7563, 23.7412, 23.7167, 23.6985, 23.6824, 23.6161, 23.5427, 23.5178, 23.4941, 23.4435, 23.3704, 23.3539, 23.3088, 23.2722, 23.2477, 23.233, 23.2335, 23.2295, 23.2211, 23.2293, 23.2299, 23.2268, 23.2175, 23.1978, 23.1826, 23.1768, 23.187, 23.1804, 23.1736, 23.115, 22.9617, 22.8332, 22.7596, 22.7407, 22.7447}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0}
}
