netcdf file-166.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (27 currently)
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391}
TIME =
  {22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556, 22579.193993055556}
TEMP =
  {25.5347, 25.5385, 25.4894, 25.4076, 25.2758, 25.1667, 25.1123, 25.0878, 25.0718, 25.0605, 25.0524, 25.0433, 25.0406, 25.0401, 25.0392, 25.0372, 25.037, 25.0367, 25.0366, 25.0366, 25.0368, 25.037, 25.0378, 25.0389, 25.0396, 25.0403, 25.0422}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.859, 23.853, 24.847, 25.841, 26.835}
}
