netcdf IMOS_ANMN-TS_20150113T230000Z_NRSROT-ADCP_FV01_NRSROT-ADCP-1409-RBR-TR-1050-43_END-20150128T062000Z_id-7741.nc {
  dimensions:
    TIME = UNLIMITED;   // (4121 currently)
  variables:
    double TIME(TIME=4121);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=4121);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=4121);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=4121);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=4121);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=4121);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=4121);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=4121);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=4121);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=4121);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=4121);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=4121);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=4121);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been filled using the DEPTH median (mooring).";
  :instrument = "RBR TR-1050";
  :references = "http://www.imos.org.au";
  :site_code = "NRSROT";
  :platform_code = "NRSROT-ADCP";
  :deployment_code = "NRSROT-ADCP-1409";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "tr20584";
  :history = "2015-01-29T09:15:56Z - depthPP: Depth computed from the only pressure sensor available, using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :geospatial_lat_min = -31.9966; // double
  :geospatial_lat_max = -31.9966; // double
  :geospatial_lon_min = 115.4157166667; // double
  :geospatial_lon_max = 115.4157166667; // double
  :instrument_nominal_depth = 43.0f; // float
  :site_nominal_depth = 48.0f; // float
  :geospatial_vertical_min = -1.338954f; // float
  :geospatial_vertical_max = 40.051956f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-09-19T05:00:00Z";
  :time_deployment_end = "2015-01-28T03:00:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-28T06:20:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.961805555555, 23753.965277777777, 23753.96875, 23753.972222222223, 23753.975694444445, 23753.979166666668, 23753.98263888889, 23753.98611111111, 23753.989583333332, 23753.993055555555, 23753.996527777777, 23754.0, 23754.003472222223, 23754.006944444445, 23754.010416666668, 23754.01388888889, 23754.01736111111, 23754.020833333332, 23754.024305555555, 23754.027777777777, 23754.03125, 23754.034722222223, 23754.038194444445, 23754.041666666668, 23754.04513888889, 23754.04861111111, 23754.052083333332, 23754.055555555555, 23754.059027777777, 23754.0625, 23754.065972222223, 23754.069444444445, 23754.072916666668, 23754.07638888889, 23754.07986111111, 23754.083333333332, 23754.086805555555, 23754.090277777777, 23754.09375, 23754.097222222223, 23754.100694444445, 23754.104166666668, 23754.10763888889, 23754.11111111111, 23754.114583333332, 23754.118055555555, 23754.121527777777, 23754.125, 23754.128472222223, 23754.131944444445, 23754.135416666668, 23754.13888888889, 23754.14236111111, 23754.145833333332, 23754.149305555555, 23754.152777777777, 23754.15625, 23754.159722222223, 23754.163194444445, 23754.166666666668, 23754.17013888889, 23754.17361111111, 23754.177083333332, 23754.180555555555, 23754.184027777777, 23754.1875, 23754.190972222223, 23754.194444444445, 23754.197916666668, 23754.20138888889, 23754.20486111111, 23754.208333333332, 23754.211805555555, 23754.215277777777, 23754.21875, 23754.222222222223, 23754.225694444445, 23754.229166666668, 23754.23263888889, 23754.23611111111, 23754.239583333332, 23754.243055555555, 23754.246527777777, 23754.25, 23754.253472222223, 23754.256944444445, 23754.260416666668, 23754.26388888889, 23754.26736111111, 23754.270833333332, 23754.274305555555, 23754.277777777777, 23754.28125, 23754.284722222223, 23754.288194444445, 23754.291666666668, 23754.29513888889, 23754.29861111111, 23754.302083333332, 23754.305555555555, 23754.309027777777, 23754.3125, 23754.315972222223, 23754.319444444445, 23754.322916666668, 23754.32638888889, 23754.32986111111, 23754.333333333332, 23754.336805555555, 23754.340277777777, 23754.34375, 23754.347222222223, 23754.350694444445, 23754.354166666668, 23754.35763888889, 23754.36111111111, 23754.364583333332, 23754.368055555555, 23754.371527777777, 23754.375, 23754.378472222223, 23754.381944444445, 23754.385416666668, 23754.38888888889, 23754.39236111111, 23754.395833333332, 23754.399305555555, 23754.402777777777, 23754.40625, 23754.409722222223, 23754.413194444445, 23754.416666666668, 23754.42013888889, 23754.42361111111, 23754.427083333332, 23754.430555555555, 23754.434027777777, 23754.4375, 23754.440972222223, 23754.444444444445, 23754.447916666668, 23754.45138888889, 23754.45486111111, 23754.458333333332, 23754.461805555555, 23754.465277777777, 23754.46875, 23754.472222222223, 23754.475694444445, 23754.479166666668, 23754.48263888889, 23754.48611111111, 23754.489583333332, 23754.493055555555, 23754.496527777777, 23754.5, 23754.503472222223, 23754.506944444445, 23754.510416666668, 23754.51388888889, 23754.51736111111, 23754.520833333332, 23754.524305555555, 23754.527777777777, 23754.53125, 23754.534722222223, 23754.538194444445, 23754.541666666668, 23754.54513888889, 23754.54861111111, 23754.552083333332, 23754.555555555555, 23754.559027777777, 23754.5625, 23754.565972222223, 23754.569444444445, 23754.572916666668, 23754.57638888889, 23754.57986111111, 23754.583333333332, 23754.586805555555, 23754.590277777777, 23754.59375, 23754.597222222223, 23754.600694444445, 23754.604166666668, 23754.60763888889, 23754.61111111111, 23754.614583333332, 23754.618055555555, 23754.621527777777, 23754.625, 23754.628472222223, 23754.631944444445, 23754.635416666668, 23754.63888888889, 23754.64236111111, 23754.645833333332, 23754.649305555555, 23754.652777777777, 23754.65625, 23754.659722222223, 23754.663194444445, 23754.666666666668, 23754.67013888889, 23754.67361111111, 23754.677083333332, 23754.680555555555, 23754.684027777777, 23754.6875, 23754.690972222223, 23754.694444444445, 23754.697916666668, 23754.70138888889, 23754.70486111111, 23754.708333333332, 23754.711805555555, 23754.715277777777, 23754.71875, 23754.722222222223, 23754.725694444445, 23754.729166666668, 23754.73263888889, 23754.73611111111, 23754.739583333332, 23754.743055555555, 23754.746527777777, 23754.75, 23754.753472222223, 23754.756944444445, 23754.760416666668, 23754.76388888889, 23754.76736111111, 23754.770833333332, 23754.774305555555, 23754.777777777777, 23754.78125, 23754.784722222223, 23754.788194444445, 23754.791666666668, 23754.79513888889, 23754.79861111111, 23754.802083333332, 23754.805555555555, 23754.809027777777, 23754.8125, 23754.815972222223, 23754.819444444445, 23754.822916666668, 23754.82638888889, 23754.82986111111, 23754.833333333332, 23754.836805555555, 23754.840277777777, 23754.84375, 23754.847222222223, 23754.850694444445, 23754.854166666668, 23754.85763888889, 23754.86111111111, 23754.864583333332, 23754.868055555555, 23754.871527777777, 23754.875, 23754.878472222223, 23754.881944444445, 23754.885416666668, 23754.88888888889, 23754.89236111111, 23754.895833333332, 23754.899305555555, 23754.902777777777, 23754.90625, 23754.909722222223, 23754.913194444445, 23754.916666666668, 23754.92013888889, 23754.92361111111, 23754.927083333332, 23754.930555555555, 23754.934027777777, 23754.9375, 23754.940972222223, 23754.944444444445, 23754.947916666668, 23754.95138888889, 23754.95486111111, 23754.958333333332, 23754.961805555555, 23754.965277777777, 23754.96875, 23754.972222222223, 23754.975694444445, 23754.979166666668, 23754.98263888889, 23754.98611111111, 23754.989583333332, 23754.993055555555, 23754.996527777777, 23755.0, 23755.003472222223, 23755.006944444445, 23755.010416666668, 23755.01388888889, 23755.01736111111, 23755.020833333332, 23755.024305555555, 23755.027777777777, 23755.03125, 23755.034722222223, 23755.038194444445, 23755.041666666668, 23755.04513888889, 23755.04861111111, 23755.052083333332, 23755.055555555555, 23755.059027777777, 23755.0625, 23755.065972222223, 23755.069444444445, 23755.072916666668, 23755.07638888889, 23755.07986111111, 23755.083333333332, 23755.086805555555, 23755.090277777777, 23755.09375, 23755.097222222223, 23755.100694444445, 23755.104166666668, 23755.10763888889, 23755.11111111111, 23755.114583333332, 23755.118055555555, 23755.121527777777, 23755.125, 23755.128472222223, 23755.131944444445, 23755.135416666668, 23755.13888888889, 23755.14236111111, 23755.145833333332, 23755.149305555555, 23755.152777777777, 23755.15625, 23755.159722222223, 23755.163194444445, 23755.166666666668, 23755.17013888889, 23755.17361111111, 23755.177083333332, 23755.180555555555, 23755.184027777777, 23755.1875, 23755.190972222223, 23755.194444444445, 23755.197916666668, 23755.20138888889, 23755.20486111111, 23755.208333333332, 23755.211805555555, 23755.215277777777, 23755.21875, 23755.222222222223, 23755.225694444445, 23755.229166666668, 23755.23263888889, 23755.23611111111, 23755.239583333332, 23755.243055555555, 23755.246527777777, 23755.25, 23755.253472222223, 23755.256944444445, 23755.260416666668, 23755.26388888889, 23755.26736111111, 23755.270833333332, 23755.274305555555, 23755.277777777777, 23755.28125, 23755.284722222223, 23755.288194444445, 23755.291666666668, 23755.29513888889, 23755.29861111111, 23755.302083333332, 23755.305555555555, 23755.309027777777, 23755.3125, 23755.315972222223, 23755.319444444445, 23755.322916666668, 23755.32638888889, 23755.32986111111, 23755.333333333332, 23755.336805555555, 23755.340277777777, 23755.34375, 23755.347222222223, 23755.350694444445, 23755.354166666668, 23755.35763888889, 23755.36111111111, 23755.364583333332, 23755.368055555555, 23755.371527777777, 23755.375, 23755.378472222223, 23755.381944444445, 23755.385416666668, 23755.38888888889, 23755.39236111111, 23755.395833333332, 23755.399305555555, 23755.402777777777, 23755.40625, 23755.409722222223, 23755.413194444445, 23755.416666666668, 23755.42013888889, 23755.42361111111, 23755.427083333332, 23755.430555555555, 23755.434027777777, 23755.4375, 23755.440972222223, 23755.444444444445, 23755.447916666668, 23755.45138888889, 23755.45486111111, 23755.458333333332, 23755.461805555555, 23755.465277777777, 23755.46875, 23755.472222222223, 23755.475694444445, 23755.479166666668, 23755.48263888889, 23755.48611111111, 23755.489583333332, 23755.493055555555, 23755.496527777777, 23755.5, 23755.503472222223, 23755.506944444445, 23755.510416666668, 23755.51388888889, 23755.51736111111, 23755.520833333332, 23755.524305555555, 23755.527777777777, 23755.53125, 23755.534722222223, 23755.538194444445, 23755.541666666668, 23755.54513888889, 23755.54861111111, 23755.552083333332, 23755.555555555555, 23755.559027777777, 23755.5625, 23755.565972222223, 23755.569444444445, 23755.572916666668, 23755.57638888889, 23755.57986111111, 23755.583333333332, 23755.586805555555, 23755.590277777777, 23755.59375, 23755.597222222223, 23755.600694444445, 23755.604166666668, 23755.60763888889, 23755.61111111111, 23755.614583333332, 23755.618055555555, 23755.621527777777, 23755.625, 23755.628472222223, 23755.631944444445, 23755.635416666668, 23755.63888888889, 23755.64236111111, 23755.645833333332, 23755.649305555555, 23755.652777777777, 23755.65625, 23755.659722222223, 23755.663194444445, 23755.666666666668, 23755.67013888889, 23755.67361111111, 23755.677083333332, 23755.680555555555, 23755.684027777777, 23755.6875, 23755.690972222223, 23755.694444444445, 23755.697916666668, 23755.70138888889, 23755.70486111111, 23755.708333333332, 23755.711805555555, 23755.715277777777, 23755.71875, 23755.722222222223, 23755.725694444445, 23755.729166666668, 23755.73263888889, 23755.73611111111, 23755.739583333332, 23755.743055555555, 23755.746527777777, 23755.75, 23755.753472222223, 23755.756944444445, 23755.760416666668, 23755.76388888889, 23755.76736111111, 23755.770833333332, 23755.774305555555, 23755.777777777777, 23755.78125, 23755.784722222223, 23755.788194444445, 23755.791666666668, 23755.79513888889, 23755.79861111111, 23755.802083333332, 23755.805555555555, 23755.809027777777, 23755.8125, 23755.815972222223, 23755.819444444445, 23755.822916666668, 23755.82638888889, 23755.82986111111, 23755.833333333332, 23755.836805555555, 23755.840277777777, 23755.84375, 23755.847222222223, 23755.850694444445, 23755.854166666668, 23755.85763888889, 23755.86111111111, 23755.864583333332, 23755.868055555555, 23755.871527777777, 23755.875, 23755.878472222223, 23755.881944444445, 23755.885416666668, 23755.88888888889, 23755.89236111111, 23755.895833333332, 23755.899305555555, 23755.902777777777, 23755.90625, 23755.909722222223, 23755.913194444445, 23755.916666666668, 23755.92013888889, 23755.92361111111, 23755.927083333332, 23755.930555555555, 23755.934027777777, 23755.9375, 23755.940972222223, 23755.944444444445, 23755.947916666668, 23755.95138888889, 23755.95486111111, 23755.958333333332, 23755.961805555555, 23755.965277777777, 23755.96875, 23755.972222222223, 23755.975694444445, 23755.979166666668, 23755.98263888889, 23755.98611111111, 23755.989583333332, 23755.993055555555, 23755.996527777777, 23756.0, 23756.003472222223, 23756.006944444445, 23756.010416666668, 23756.01388888889, 23756.01736111111, 23756.020833333332, 23756.024305555555, 23756.027777777777, 23756.03125, 23756.034722222223, 23756.038194444445, 23756.041666666668, 23756.04513888889, 23756.04861111111, 23756.052083333332, 23756.055555555555, 23756.059027777777, 23756.0625, 23756.065972222223, 23756.069444444445, 23756.072916666668, 23756.07638888889, 23756.07986111111, 23756.083333333332, 23756.086805555555, 23756.090277777777, 23756.09375, 23756.097222222223, 23756.100694444445, 23756.104166666668, 23756.10763888889, 23756.11111111111, 23756.114583333332, 23756.118055555555, 23756.121527777777, 23756.125, 23756.128472222223, 23756.131944444445, 23756.135416666668, 23756.13888888889, 23756.14236111111, 23756.145833333332, 23756.149305555555, 23756.152777777777, 23756.15625, 23756.159722222223, 23756.163194444445, 23756.166666666668, 23756.17013888889, 23756.17361111111, 23756.177083333332, 23756.180555555555, 23756.184027777777, 23756.1875, 23756.190972222223, 23756.194444444445, 23756.197916666668, 23756.20138888889, 23756.20486111111, 23756.208333333332, 23756.211805555555, 23756.215277777777, 23756.21875, 23756.222222222223, 23756.225694444445, 23756.229166666668, 23756.23263888889, 23756.23611111111, 23756.239583333332, 23756.243055555555, 23756.246527777777, 23756.25, 23756.253472222223, 23756.256944444445, 23756.260416666668, 23756.26388888889, 23756.26736111111, 23756.270833333332, 23756.274305555555, 23756.277777777777, 23756.28125, 23756.284722222223, 23756.288194444445, 23756.291666666668, 23756.29513888889, 23756.29861111111, 23756.302083333332, 23756.305555555555, 23756.309027777777, 23756.3125, 23756.315972222223, 23756.319444444445, 23756.322916666668, 23756.32638888889, 23756.32986111111, 23756.333333333332, 23756.336805555555, 23756.340277777777, 23756.34375, 23756.347222222223, 23756.350694444445, 23756.354166666668, 23756.35763888889, 23756.36111111111, 23756.364583333332, 23756.368055555555, 23756.371527777777, 23756.375, 23756.378472222223, 23756.381944444445, 23756.385416666668, 23756.38888888889, 23756.39236111111, 23756.395833333332, 23756.399305555555, 23756.402777777777, 23756.40625, 23756.409722222223, 23756.413194444445, 23756.416666666668, 23756.42013888889, 23756.42361111111, 23756.427083333332, 23756.430555555555, 23756.434027777777, 23756.4375, 23756.440972222223, 23756.444444444445, 23756.447916666668, 23756.45138888889, 23756.45486111111, 23756.458333333332, 23756.461805555555, 23756.465277777777, 23756.46875, 23756.472222222223, 23756.475694444445, 23756.479166666668, 23756.48263888889, 23756.48611111111, 23756.489583333332, 23756.493055555555, 23756.496527777777, 23756.5, 23756.503472222223, 23756.506944444445, 23756.510416666668, 23756.51388888889, 23756.51736111111, 23756.520833333332, 23756.524305555555, 23756.527777777777, 23756.53125, 23756.534722222223, 23756.538194444445, 23756.541666666668, 23756.54513888889, 23756.54861111111, 23756.552083333332, 23756.555555555555, 23756.559027777777, 23756.5625, 23756.565972222223, 23756.569444444445, 23756.572916666668, 23756.57638888889, 23756.57986111111, 23756.583333333332, 23756.586805555555, 23756.590277777777, 23756.59375, 23756.597222222223, 23756.600694444445, 23756.604166666668, 23756.60763888889, 23756.61111111111, 23756.614583333332, 23756.618055555555, 23756.621527777777, 23756.625, 23756.628472222223, 23756.631944444445, 23756.635416666668, 23756.63888888889, 23756.64236111111, 23756.645833333332, 23756.649305555555, 23756.652777777777, 23756.65625, 23756.659722222223, 23756.663194444445, 23756.666666666668, 23756.67013888889, 23756.67361111111, 23756.677083333332, 23756.680555555555, 23756.684027777777, 23756.6875, 23756.690972222223, 23756.694444444445, 23756.697916666668, 23756.70138888889, 23756.70486111111, 23756.708333333332, 23756.711805555555, 23756.715277777777, 23756.71875, 23756.722222222223, 23756.725694444445, 23756.729166666668, 23756.73263888889, 23756.73611111111, 23756.739583333332, 23756.743055555555, 23756.746527777777, 23756.75, 23756.753472222223, 23756.756944444445, 23756.760416666668, 23756.76388888889, 23756.76736111111, 23756.770833333332, 23756.774305555555, 23756.777777777777, 23756.78125, 23756.784722222223, 23756.788194444445, 23756.791666666668, 23756.79513888889, 23756.79861111111, 23756.802083333332, 23756.805555555555, 23756.809027777777, 23756.8125, 23756.815972222223, 23756.819444444445, 23756.822916666668, 23756.82638888889, 23756.82986111111, 23756.833333333332, 23756.836805555555, 23756.840277777777, 23756.84375, 23756.847222222223, 23756.850694444445, 23756.854166666668, 23756.85763888889, 23756.86111111111, 23756.864583333332, 23756.868055555555, 23756.871527777777, 23756.875, 23756.878472222223, 23756.881944444445, 23756.885416666668, 23756.88888888889, 23756.89236111111, 23756.895833333332, 23756.899305555555, 23756.902777777777, 23756.90625, 23756.909722222223, 23756.913194444445, 23756.916666666668, 23756.92013888889, 23756.92361111111, 23756.927083333332, 23756.930555555555, 23756.934027777777, 23756.9375, 23756.940972222223, 23756.944444444445, 23756.947916666668, 23756.95138888889, 23756.95486111111, 23756.958333333332, 23756.961805555555, 23756.965277777777, 23756.96875, 23756.972222222223, 23756.975694444445, 23756.979166666668, 23756.98263888889, 23756.98611111111, 23756.989583333332, 23756.993055555555, 23756.996527777777, 23757.0, 23757.003472222223, 23757.006944444445, 23757.010416666668, 23757.01388888889, 23757.01736111111, 23757.020833333332, 23757.024305555555, 23757.027777777777, 23757.03125, 23757.034722222223, 23757.038194444445, 23757.041666666668, 23757.04513888889, 23757.04861111111, 23757.052083333332, 23757.055555555555, 23757.059027777777, 23757.0625, 23757.065972222223, 23757.069444444445, 23757.072916666668, 23757.07638888889, 23757.07986111111, 23757.083333333332, 23757.086805555555, 23757.090277777777, 23757.09375, 23757.097222222223, 23757.100694444445, 23757.104166666668, 23757.10763888889, 23757.11111111111, 23757.114583333332, 23757.118055555555, 23757.121527777777, 23757.125, 23757.128472222223, 23757.131944444445, 23757.135416666668, 23757.13888888889, 23757.14236111111, 23757.145833333332, 23757.149305555555, 23757.152777777777, 23757.15625, 23757.159722222223, 23757.163194444445, 23757.166666666668, 23757.17013888889, 23757.17361111111, 23757.177083333332, 23757.180555555555, 23757.184027777777, 23757.1875, 23757.190972222223, 23757.194444444445, 23757.197916666668, 23757.20138888889, 23757.20486111111, 23757.208333333332, 23757.211805555555, 23757.215277777777, 23757.21875, 23757.222222222223, 23757.225694444445, 23757.229166666668, 23757.23263888889, 23757.23611111111, 23757.239583333332, 23757.243055555555, 23757.246527777777, 23757.25, 23757.253472222223, 23757.256944444445, 23757.260416666668, 23757.26388888889, 23757.26736111111, 23757.270833333332, 23757.274305555555, 23757.277777777777, 23757.28125, 23757.284722222223, 23757.288194444445, 23757.291666666668, 23757.29513888889, 23757.29861111111, 23757.302083333332, 23757.305555555555, 23757.309027777777, 23757.3125, 23757.315972222223, 23757.319444444445, 23757.322916666668, 23757.32638888889, 23757.32986111111, 23757.333333333332, 23757.336805555555, 23757.340277777777, 23757.34375, 23757.347222222223, 23757.350694444445, 23757.354166666668, 23757.35763888889, 23757.36111111111, 23757.364583333332, 23757.368055555555, 23757.371527777777, 23757.375, 23757.378472222223, 23757.381944444445, 23757.385416666668, 23757.38888888889, 23757.39236111111, 23757.395833333332, 23757.399305555555, 23757.402777777777, 23757.40625, 23757.409722222223, 23757.413194444445, 23757.416666666668, 23757.42013888889, 23757.42361111111, 23757.427083333332, 23757.430555555555, 23757.434027777777, 23757.4375, 23757.440972222223, 23757.444444444445, 23757.447916666668, 23757.45138888889, 23757.45486111111, 23757.458333333332, 23757.461805555555, 23757.465277777777, 23757.46875, 23757.472222222223, 23757.475694444445, 23757.479166666668, 23757.48263888889, 23757.48611111111, 23757.489583333332, 23757.493055555555, 23757.496527777777, 23757.5, 23757.503472222223, 23757.506944444445, 23757.510416666668, 23757.51388888889, 23757.51736111111, 23757.520833333332, 23757.524305555555, 23757.527777777777, 23757.53125, 23757.534722222223, 23757.538194444445, 23757.541666666668, 23757.54513888889, 23757.54861111111, 23757.552083333332, 23757.555555555555, 23757.559027777777, 23757.5625, 23757.565972222223, 23757.569444444445, 23757.572916666668, 23757.57638888889, 23757.57986111111, 23757.583333333332, 23757.586805555555, 23757.590277777777, 23757.59375, 23757.597222222223, 23757.600694444445, 23757.604166666668, 23757.60763888889, 23757.61111111111, 23757.614583333332, 23757.618055555555, 23757.621527777777, 23757.625, 23757.628472222223, 23757.631944444445, 23757.635416666668, 23757.63888888889, 23757.64236111111, 23757.645833333332, 23757.649305555555, 23757.652777777777, 23757.65625, 23757.659722222223, 23757.663194444445, 23757.666666666668, 23757.67013888889, 23757.67361111111, 23757.677083333332, 23757.680555555555, 23757.684027777777, 23757.6875, 23757.690972222223, 23757.694444444445, 23757.697916666668, 23757.70138888889, 23757.70486111111, 23757.708333333332, 23757.711805555555, 23757.715277777777, 23757.71875, 23757.722222222223, 23757.725694444445, 23757.729166666668, 23757.73263888889, 23757.73611111111, 23757.739583333332, 23757.743055555555, 23757.746527777777, 23757.75, 23757.753472222223, 23757.756944444445, 23757.760416666668, 23757.76388888889, 23757.76736111111, 23757.770833333332, 23757.774305555555, 23757.777777777777, 23757.78125, 23757.784722222223, 23757.788194444445, 23757.791666666668, 23757.79513888889, 23757.79861111111, 23757.802083333332, 23757.805555555555, 23757.809027777777, 23757.8125, 23757.815972222223, 23757.819444444445, 23757.822916666668, 23757.82638888889, 23757.82986111111, 23757.833333333332, 23757.836805555555, 23757.840277777777, 23757.84375, 23757.847222222223, 23757.850694444445, 23757.854166666668, 23757.85763888889, 23757.86111111111, 23757.864583333332, 23757.868055555555, 23757.871527777777, 23757.875, 23757.878472222223, 23757.881944444445, 23757.885416666668, 23757.88888888889, 23757.89236111111, 23757.895833333332, 23757.899305555555, 23757.902777777777, 23757.90625, 23757.909722222223, 23757.913194444445, 23757.916666666668, 23757.92013888889, 23757.92361111111, 23757.927083333332, 23757.930555555555, 23757.934027777777, 23757.9375, 23757.940972222223, 23757.944444444445, 23757.947916666668, 23757.95138888889, 23757.95486111111, 23757.958333333332, 23757.961805555555, 23757.965277777777, 23757.96875, 23757.972222222223, 23757.975694444445, 23757.979166666668, 23757.98263888889, 23757.98611111111, 23757.989583333332, 23757.993055555555, 23757.996527777777, 23758.0, 23758.003472222223, 23758.006944444445, 23758.010416666668, 23758.01388888889, 23758.01736111111, 23758.020833333332, 23758.024305555555, 23758.027777777777, 23758.03125, 23758.034722222223, 23758.038194444445, 23758.041666666668, 23758.04513888889, 23758.04861111111, 23758.052083333332, 23758.055555555555, 23758.059027777777, 23758.0625, 23758.065972222223, 23758.069444444445, 23758.072916666668, 23758.07638888889, 23758.07986111111, 23758.083333333332, 23758.086805555555, 23758.090277777777, 23758.09375, 23758.097222222223, 23758.100694444445, 23758.104166666668, 23758.10763888889, 23758.11111111111, 23758.114583333332, 23758.118055555555, 23758.121527777777, 23758.125, 23758.128472222223, 23758.131944444445, 23758.135416666668, 23758.13888888889, 23758.14236111111, 23758.145833333332, 23758.149305555555, 23758.152777777777, 23758.15625, 23758.159722222223, 23758.163194444445, 23758.166666666668, 23758.17013888889, 23758.17361111111, 23758.177083333332, 23758.180555555555, 23758.184027777777, 23758.1875, 23758.190972222223, 23758.194444444445, 23758.197916666668, 23758.20138888889, 23758.20486111111, 23758.208333333332, 23758.211805555555, 23758.215277777777, 23758.21875, 23758.222222222223, 23758.225694444445, 23758.229166666668, 23758.23263888889, 23758.23611111111, 23758.239583333332, 23758.243055555555, 23758.246527777777, 23758.25, 23758.253472222223, 23758.256944444445, 23758.260416666668, 23758.26388888889, 23758.26736111111, 23758.270833333332, 23758.274305555555, 23758.277777777777, 23758.28125, 23758.284722222223, 23758.288194444445, 23758.291666666668, 23758.29513888889, 23758.29861111111, 23758.302083333332, 23758.305555555555, 23758.309027777777, 23758.3125, 23758.315972222223, 23758.319444444445, 23758.322916666668, 23758.32638888889, 23758.32986111111, 23758.333333333332, 23758.336805555555, 23758.340277777777, 23758.34375, 23758.347222222223, 23758.350694444445, 23758.354166666668, 23758.35763888889, 23758.36111111111, 23758.364583333332, 23758.368055555555, 23758.371527777777, 23758.375, 23758.378472222223, 23758.381944444445, 23758.385416666668, 23758.38888888889, 23758.39236111111, 23758.395833333332, 23758.399305555555, 23758.402777777777, 23758.40625, 23758.409722222223, 23758.413194444445, 23758.416666666668, 23758.42013888889, 23758.42361111111, 23758.427083333332, 23758.430555555555, 23758.434027777777, 23758.4375, 23758.440972222223, 23758.444444444445, 23758.447916666668, 23758.45138888889, 23758.45486111111, 23758.458333333332, 23758.461805555555, 23758.465277777777, 23758.46875, 23758.472222222223, 23758.475694444445, 23758.479166666668, 23758.48263888889, 23758.48611111111, 23758.489583333332, 23758.493055555555, 23758.496527777777, 23758.5, 23758.503472222223, 23758.506944444445, 23758.510416666668, 23758.51388888889, 23758.51736111111, 23758.520833333332, 23758.524305555555, 23758.527777777777, 23758.53125, 23758.534722222223, 23758.538194444445, 23758.541666666668, 23758.54513888889, 23758.54861111111, 23758.552083333332, 23758.555555555555, 23758.559027777777, 23758.5625, 23758.565972222223, 23758.569444444445, 23758.572916666668, 23758.57638888889, 23758.57986111111, 23758.583333333332, 23758.586805555555, 23758.590277777777, 23758.59375, 23758.597222222223, 23758.600694444445, 23758.604166666668, 23758.60763888889, 23758.61111111111, 23758.614583333332, 23758.618055555555, 23758.621527777777, 23758.625, 23758.628472222223, 23758.631944444445, 23758.635416666668, 23758.63888888889, 23758.64236111111, 23758.645833333332, 23758.649305555555, 23758.652777777777, 23758.65625, 23758.659722222223, 23758.663194444445, 23758.666666666668, 23758.67013888889, 23758.67361111111, 23758.677083333332, 23758.680555555555, 23758.684027777777, 23758.6875, 23758.690972222223, 23758.694444444445, 23758.697916666668, 23758.70138888889, 23758.70486111111, 23758.708333333332, 23758.711805555555, 23758.715277777777, 23758.71875, 23758.722222222223, 23758.725694444445, 23758.729166666668, 23758.73263888889, 23758.73611111111, 23758.739583333332, 23758.743055555555, 23758.746527777777, 23758.75, 23758.753472222223, 23758.756944444445, 23758.760416666668, 23758.76388888889, 23758.76736111111, 23758.770833333332, 23758.774305555555, 23758.777777777777, 23758.78125, 23758.784722222223, 23758.788194444445, 23758.791666666668, 23758.79513888889, 23758.79861111111, 23758.802083333332, 23758.805555555555, 23758.809027777777, 23758.8125, 23758.815972222223, 23758.819444444445, 23758.822916666668, 23758.82638888889, 23758.82986111111, 23758.833333333332, 23758.836805555555, 23758.840277777777, 23758.84375, 23758.847222222223, 23758.850694444445, 23758.854166666668, 23758.85763888889, 23758.86111111111, 23758.864583333332, 23758.868055555555, 23758.871527777777, 23758.875, 23758.878472222223, 23758.881944444445, 23758.885416666668, 23758.88888888889, 23758.89236111111, 23758.895833333332, 23758.899305555555, 23758.902777777777, 23758.90625, 23758.909722222223, 23758.913194444445, 23758.916666666668, 23758.92013888889, 23758.92361111111, 23758.927083333332, 23758.930555555555, 23758.934027777777, 23758.9375, 23758.940972222223, 23758.944444444445, 23758.947916666668, 23758.95138888889, 23758.95486111111, 23758.958333333332, 23758.961805555555, 23758.965277777777, 23758.96875, 23758.972222222223, 23758.975694444445, 23758.979166666668, 23758.98263888889, 23758.98611111111, 23758.989583333332, 23758.993055555555, 23758.996527777777, 23759.0, 23759.003472222223, 23759.006944444445, 23759.010416666668, 23759.01388888889, 23759.01736111111, 23759.020833333332, 23759.024305555555, 23759.027777777777, 23759.03125, 23759.034722222223, 23759.038194444445, 23759.041666666668, 23759.04513888889, 23759.04861111111, 23759.052083333332, 23759.055555555555, 23759.059027777777, 23759.0625, 23759.065972222223, 23759.069444444445, 23759.072916666668, 23759.07638888889, 23759.07986111111, 23759.083333333332, 23759.086805555555, 23759.090277777777, 23759.09375, 23759.097222222223, 23759.100694444445, 23759.104166666668, 23759.10763888889, 23759.11111111111, 23759.114583333332, 23759.118055555555, 23759.121527777777, 23759.125, 23759.128472222223, 23759.131944444445, 23759.135416666668, 23759.13888888889, 23759.14236111111, 23759.145833333332, 23759.149305555555, 23759.152777777777, 23759.15625, 23759.159722222223, 23759.163194444445, 23759.166666666668, 23759.17013888889, 23759.17361111111, 23759.177083333332, 23759.180555555555, 23759.184027777777, 23759.1875, 23759.190972222223, 23759.194444444445, 23759.197916666668, 23759.20138888889, 23759.20486111111, 23759.208333333332, 23759.211805555555, 23759.215277777777, 23759.21875, 23759.222222222223, 23759.225694444445, 23759.229166666668, 23759.23263888889, 23759.23611111111, 23759.239583333332, 23759.243055555555, 23759.246527777777, 23759.25, 23759.253472222223, 23759.256944444445, 23759.260416666668, 23759.26388888889, 23759.26736111111, 23759.270833333332, 23759.274305555555, 23759.277777777777, 23759.28125, 23759.284722222223, 23759.288194444445, 23759.291666666668, 23759.29513888889, 23759.29861111111, 23759.302083333332, 23759.305555555555, 23759.309027777777, 23759.3125, 23759.315972222223, 23759.319444444445, 23759.322916666668, 23759.32638888889, 23759.32986111111, 23759.333333333332, 23759.336805555555, 23759.340277777777, 23759.34375, 23759.347222222223, 23759.350694444445, 23759.354166666668, 23759.35763888889, 23759.36111111111, 23759.364583333332, 23759.368055555555, 23759.371527777777, 23759.375, 23759.378472222223, 23759.381944444445, 23759.385416666668, 23759.38888888889, 23759.39236111111, 23759.395833333332, 23759.399305555555, 23759.402777777777, 23759.40625, 23759.409722222223, 23759.413194444445, 23759.416666666668, 23759.42013888889, 23759.42361111111, 23759.427083333332, 23759.430555555555, 23759.434027777777, 23759.4375, 23759.440972222223, 23759.444444444445, 23759.447916666668, 23759.45138888889, 23759.45486111111, 23759.458333333332, 23759.461805555555, 23759.465277777777, 23759.46875, 23759.472222222223, 23759.475694444445, 23759.479166666668, 23759.48263888889, 23759.48611111111, 23759.489583333332, 23759.493055555555, 23759.496527777777, 23759.5, 23759.503472222223, 23759.506944444445, 23759.510416666668, 23759.51388888889, 23759.51736111111, 23759.520833333332, 23759.524305555555, 23759.527777777777, 23759.53125, 23759.534722222223, 23759.538194444445, 23759.541666666668, 23759.54513888889, 23759.54861111111, 23759.552083333332, 23759.555555555555, 23759.559027777777, 23759.5625, 23759.565972222223, 23759.569444444445, 23759.572916666668, 23759.57638888889, 23759.57986111111, 23759.583333333332, 23759.586805555555, 23759.590277777777, 23759.59375, 23759.597222222223, 23759.600694444445, 23759.604166666668, 23759.60763888889, 23759.61111111111, 23759.614583333332, 23759.618055555555, 23759.621527777777, 23759.625, 23759.628472222223, 23759.631944444445, 23759.635416666668, 23759.63888888889, 23759.64236111111, 23759.645833333332, 23759.649305555555, 23759.652777777777, 23759.65625, 23759.659722222223, 23759.663194444445, 23759.666666666668, 23759.67013888889, 23759.67361111111, 23759.677083333332, 23759.680555555555, 23759.684027777777, 23759.6875, 23759.690972222223, 23759.694444444445, 23759.697916666668, 23759.70138888889, 23759.70486111111, 23759.708333333332, 23759.711805555555, 23759.715277777777, 23759.71875, 23759.722222222223, 23759.725694444445, 23759.729166666668, 23759.73263888889, 23759.73611111111, 23759.739583333332, 23759.743055555555, 23759.746527777777, 23759.75, 23759.753472222223, 23759.756944444445, 23759.760416666668, 23759.76388888889, 23759.76736111111, 23759.770833333332, 23759.774305555555, 23759.777777777777, 23759.78125, 23759.784722222223, 23759.788194444445, 23759.791666666668, 23759.79513888889, 23759.79861111111, 23759.802083333332, 23759.805555555555, 23759.809027777777, 23759.8125, 23759.815972222223, 23759.819444444445, 23759.822916666668, 23759.82638888889, 23759.82986111111, 23759.833333333332, 23759.836805555555, 23759.840277777777, 23759.84375, 23759.847222222223, 23759.850694444445, 23759.854166666668, 23759.85763888889, 23759.86111111111, 23759.864583333332, 23759.868055555555, 23759.871527777777, 23759.875, 23759.878472222223, 23759.881944444445, 23759.885416666668, 23759.88888888889, 23759.89236111111, 23759.895833333332, 23759.899305555555, 23759.902777777777, 23759.90625, 23759.909722222223, 23759.913194444445, 23759.916666666668, 23759.92013888889, 23759.92361111111, 23759.927083333332, 23759.930555555555, 23759.934027777777, 23759.9375, 23759.940972222223, 23759.944444444445, 23759.947916666668, 23759.95138888889, 23759.95486111111, 23759.958333333332, 23759.961805555555, 23759.965277777777, 23759.96875, 23759.972222222223, 23759.975694444445, 23759.979166666668, 23759.98263888889, 23759.98611111111, 23759.989583333332, 23759.993055555555, 23759.996527777777, 23760.0, 23760.003472222223, 23760.006944444445, 23760.010416666668, 23760.01388888889, 23760.01736111111, 23760.020833333332, 23760.024305555555, 23760.027777777777, 23760.03125, 23760.034722222223, 23760.038194444445, 23760.041666666668, 23760.04513888889, 23760.04861111111, 23760.052083333332, 23760.055555555555, 23760.059027777777, 23760.0625, 23760.065972222223, 23760.069444444445, 23760.072916666668, 23760.07638888889, 23760.07986111111, 23760.083333333332, 23760.086805555555, 23760.090277777777, 23760.09375, 23760.097222222223, 23760.100694444445, 23760.104166666668, 23760.10763888889, 23760.11111111111, 23760.114583333332, 23760.118055555555, 23760.121527777777, 23760.125, 23760.128472222223, 23760.131944444445, 23760.135416666668, 23760.13888888889, 23760.14236111111, 23760.145833333332, 23760.149305555555, 23760.152777777777, 23760.15625, 23760.159722222223, 23760.163194444445, 23760.166666666668, 23760.17013888889, 23760.17361111111, 23760.177083333332, 23760.180555555555, 23760.184027777777, 23760.1875, 23760.190972222223, 23760.194444444445, 23760.197916666668, 23760.20138888889, 23760.20486111111, 23760.208333333332, 23760.211805555555, 23760.215277777777, 23760.21875, 23760.222222222223, 23760.225694444445, 23760.229166666668, 23760.23263888889, 23760.23611111111, 23760.239583333332, 23760.243055555555, 23760.246527777777, 23760.25, 23760.253472222223, 23760.256944444445, 23760.260416666668, 23760.26388888889, 23760.26736111111, 23760.270833333332, 23760.274305555555, 23760.277777777777, 23760.28125, 23760.284722222223, 23760.288194444445, 23760.291666666668, 23760.29513888889, 23760.29861111111, 23760.302083333332, 23760.305555555555, 23760.309027777777, 23760.3125, 23760.315972222223, 23760.319444444445, 23760.322916666668, 23760.32638888889, 23760.32986111111, 23760.333333333332, 23760.336805555555, 23760.340277777777, 23760.34375, 23760.347222222223, 23760.350694444445, 23760.354166666668, 23760.35763888889, 23760.36111111111, 23760.364583333332, 23760.368055555555, 23760.371527777777, 23760.375, 23760.378472222223, 23760.381944444445, 23760.385416666668, 23760.38888888889, 23760.39236111111, 23760.395833333332, 23760.399305555555, 23760.402777777777, 23760.40625, 23760.409722222223, 23760.413194444445, 23760.416666666668, 23760.42013888889, 23760.42361111111, 23760.427083333332, 23760.430555555555, 23760.434027777777, 23760.4375, 23760.440972222223, 23760.444444444445, 23760.447916666668, 23760.45138888889, 23760.45486111111, 23760.458333333332, 23760.461805555555, 23760.465277777777, 23760.46875, 23760.472222222223, 23760.475694444445, 23760.479166666668, 23760.48263888889, 23760.48611111111, 23760.489583333332, 23760.493055555555, 23760.496527777777, 23760.5, 23760.503472222223, 23760.506944444445, 23760.510416666668, 23760.51388888889, 23760.51736111111, 23760.520833333332, 23760.524305555555, 23760.527777777777, 23760.53125, 23760.534722222223, 23760.538194444445, 23760.541666666668, 23760.54513888889, 23760.54861111111, 23760.552083333332, 23760.555555555555, 23760.559027777777, 23760.5625, 23760.565972222223, 23760.569444444445, 23760.572916666668, 23760.57638888889, 23760.57986111111, 23760.583333333332, 23760.586805555555, 23760.590277777777, 23760.59375, 23760.597222222223, 23760.600694444445, 23760.604166666668, 23760.60763888889, 23760.61111111111, 23760.614583333332, 23760.618055555555, 23760.621527777777, 23760.625, 23760.628472222223, 23760.631944444445, 23760.635416666668, 23760.63888888889, 23760.64236111111, 23760.645833333332, 23760.649305555555, 23760.652777777777, 23760.65625, 23760.659722222223, 23760.663194444445, 23760.666666666668, 23760.67013888889, 23760.67361111111, 23760.677083333332, 23760.680555555555, 23760.684027777777, 23760.6875, 23760.690972222223, 23760.694444444445, 23760.697916666668, 23760.70138888889, 23760.70486111111, 23760.708333333332, 23760.711805555555, 23760.715277777777, 23760.71875, 23760.722222222223, 23760.725694444445, 23760.729166666668, 23760.73263888889, 23760.73611111111, 23760.739583333332, 23760.743055555555, 23760.746527777777, 23760.75, 23760.753472222223, 23760.756944444445, 23760.760416666668, 23760.76388888889, 23760.76736111111, 23760.770833333332, 23760.774305555555, 23760.777777777777, 23760.78125, 23760.784722222223, 23760.788194444445, 23760.791666666668, 23760.79513888889, 23760.79861111111, 23760.802083333332, 23760.805555555555, 23760.809027777777, 23760.8125, 23760.815972222223, 23760.819444444445, 23760.822916666668, 23760.82638888889, 23760.82986111111, 23760.833333333332, 23760.836805555555, 23760.840277777777, 23760.84375, 23760.847222222223, 23760.850694444445, 23760.854166666668, 23760.85763888889, 23760.86111111111, 23760.864583333332, 23760.868055555555, 23760.871527777777, 23760.875, 23760.878472222223, 23760.881944444445, 23760.885416666668, 23760.88888888889, 23760.89236111111, 23760.895833333332, 23760.899305555555, 23760.902777777777, 23760.90625, 23760.909722222223, 23760.913194444445, 23760.916666666668, 23760.92013888889, 23760.92361111111, 23760.927083333332, 23760.930555555555, 23760.934027777777, 23760.9375, 23760.940972222223, 23760.944444444445, 23760.947916666668, 23760.95138888889, 23760.95486111111, 23760.958333333332, 23760.961805555555, 23760.965277777777, 23760.96875, 23760.972222222223, 23760.975694444445, 23760.979166666668, 23760.98263888889, 23760.98611111111, 23760.989583333332, 23760.993055555555, 23760.996527777777, 23761.0, 23761.003472222223, 23761.006944444445, 23761.010416666668, 23761.01388888889, 23761.01736111111, 23761.020833333332, 23761.024305555555, 23761.027777777777, 23761.03125, 23761.034722222223, 23761.038194444445, 23761.041666666668, 23761.04513888889, 23761.04861111111, 23761.052083333332, 23761.055555555555, 23761.059027777777, 23761.0625, 23761.065972222223, 23761.069444444445, 23761.072916666668, 23761.07638888889, 23761.07986111111, 23761.083333333332, 23761.086805555555, 23761.090277777777, 23761.09375, 23761.097222222223, 23761.100694444445, 23761.104166666668, 23761.10763888889, 23761.11111111111, 23761.114583333332, 23761.118055555555, 23761.121527777777, 23761.125, 23761.128472222223, 23761.131944444445, 23761.135416666668, 23761.13888888889, 23761.14236111111, 23761.145833333332, 23761.149305555555, 23761.152777777777, 23761.15625, 23761.159722222223, 23761.163194444445, 23761.166666666668, 23761.17013888889, 23761.17361111111, 23761.177083333332, 23761.180555555555, 23761.184027777777, 23761.1875, 23761.190972222223, 23761.194444444445, 23761.197916666668, 23761.20138888889, 23761.20486111111, 23761.208333333332, 23761.211805555555, 23761.215277777777, 23761.21875, 23761.222222222223, 23761.225694444445, 23761.229166666668, 23761.23263888889, 23761.23611111111, 23761.239583333332, 23761.243055555555, 23761.246527777777, 23761.25, 23761.253472222223, 23761.256944444445, 23761.260416666668, 23761.26388888889, 23761.26736111111, 23761.270833333332, 23761.274305555555, 23761.277777777777, 23761.28125, 23761.284722222223, 23761.288194444445, 23761.291666666668, 23761.29513888889, 23761.29861111111, 23761.302083333332, 23761.305555555555, 23761.309027777777, 23761.3125, 23761.315972222223, 23761.319444444445, 23761.322916666668, 23761.32638888889, 23761.32986111111, 23761.333333333332, 23761.336805555555, 23761.340277777777, 23761.34375, 23761.347222222223, 23761.350694444445, 23761.354166666668, 23761.35763888889, 23761.36111111111, 23761.364583333332, 23761.368055555555, 23761.371527777777, 23761.375, 23761.378472222223, 23761.381944444445, 23761.385416666668, 23761.38888888889, 23761.39236111111, 23761.395833333332, 23761.399305555555, 23761.402777777777, 23761.40625, 23761.409722222223, 23761.413194444445, 23761.416666666668, 23761.42013888889, 23761.42361111111, 23761.427083333332, 23761.430555555555, 23761.434027777777, 23761.4375, 23761.440972222223, 23761.444444444445, 23761.447916666668, 23761.45138888889, 23761.45486111111, 23761.458333333332, 23761.461805555555, 23761.465277777777, 23761.46875, 23761.472222222223, 23761.475694444445, 23761.479166666668, 23761.48263888889, 23761.48611111111, 23761.489583333332, 23761.493055555555, 23761.496527777777, 23761.5, 23761.503472222223, 23761.506944444445, 23761.510416666668, 23761.51388888889, 23761.51736111111, 23761.520833333332, 23761.524305555555, 23761.527777777777, 23761.53125, 23761.534722222223, 23761.538194444445, 23761.541666666668, 23761.54513888889, 23761.54861111111, 23761.552083333332, 23761.555555555555, 23761.559027777777, 23761.5625, 23761.565972222223, 23761.569444444445, 23761.572916666668, 23761.57638888889, 23761.57986111111, 23761.583333333332, 23761.586805555555, 23761.590277777777, 23761.59375, 23761.597222222223, 23761.600694444445, 23761.604166666668, 23761.60763888889, 23761.61111111111, 23761.614583333332, 23761.618055555555, 23761.621527777777, 23761.625, 23761.628472222223, 23761.631944444445, 23761.635416666668, 23761.63888888889, 23761.64236111111, 23761.645833333332, 23761.649305555555, 23761.652777777777, 23761.65625, 23761.659722222223, 23761.663194444445, 23761.666666666668, 23761.67013888889, 23761.67361111111, 23761.677083333332, 23761.680555555555, 23761.684027777777, 23761.6875, 23761.690972222223, 23761.694444444445, 23761.697916666668, 23761.70138888889, 23761.70486111111, 23761.708333333332, 23761.711805555555, 23761.715277777777, 23761.71875, 23761.722222222223, 23761.725694444445, 23761.729166666668, 23761.73263888889, 23761.73611111111, 23761.739583333332, 23761.743055555555, 23761.746527777777, 23761.75, 23761.753472222223, 23761.756944444445, 23761.760416666668, 23761.76388888889, 23761.76736111111, 23761.770833333332, 23761.774305555555, 23761.777777777777, 23761.78125, 23761.784722222223, 23761.788194444445, 23761.791666666668, 23761.79513888889, 23761.79861111111, 23761.802083333332, 23761.805555555555, 23761.809027777777, 23761.8125, 23761.815972222223, 23761.819444444445, 23761.822916666668, 23761.82638888889, 23761.82986111111, 23761.833333333332, 23761.836805555555, 23761.840277777777, 23761.84375, 23761.847222222223, 23761.850694444445, 23761.854166666668, 23761.85763888889, 23761.86111111111, 23761.864583333332, 23761.868055555555, 23761.871527777777, 23761.875, 23761.878472222223, 23761.881944444445, 23761.885416666668, 23761.88888888889, 23761.89236111111, 23761.895833333332, 23761.899305555555, 23761.902777777777, 23761.90625, 23761.909722222223, 23761.913194444445, 23761.916666666668, 23761.92013888889, 23761.92361111111, 23761.927083333332, 23761.930555555555, 23761.934027777777, 23761.9375, 23761.940972222223, 23761.944444444445, 23761.947916666668, 23761.95138888889, 23761.95486111111, 23761.958333333332, 23761.961805555555, 23761.965277777777, 23761.96875, 23761.972222222223, 23761.975694444445, 23761.979166666668, 23761.98263888889, 23761.98611111111, 23761.989583333332, 23761.993055555555, 23761.996527777777, 23762.0, 23762.003472222223, 23762.006944444445, 23762.010416666668, 23762.01388888889, 23762.01736111111, 23762.020833333332, 23762.024305555555, 23762.027777777777, 23762.03125, 23762.034722222223, 23762.038194444445, 23762.041666666668, 23762.04513888889, 23762.04861111111, 23762.052083333332, 23762.055555555555, 23762.059027777777, 23762.0625, 23762.065972222223, 23762.069444444445, 23762.072916666668, 23762.07638888889, 23762.07986111111, 23762.083333333332, 23762.086805555555, 23762.090277777777, 23762.09375, 23762.097222222223, 23762.100694444445, 23762.104166666668, 23762.10763888889, 23762.11111111111, 23762.114583333332, 23762.118055555555, 23762.121527777777, 23762.125, 23762.128472222223, 23762.131944444445, 23762.135416666668, 23762.13888888889, 23762.14236111111, 23762.145833333332, 23762.149305555555, 23762.152777777777, 23762.15625, 23762.159722222223, 23762.163194444445, 23762.166666666668, 23762.17013888889, 23762.17361111111, 23762.177083333332, 23762.180555555555, 23762.184027777777, 23762.1875, 23762.190972222223, 23762.194444444445, 23762.197916666668, 23762.20138888889, 23762.20486111111, 23762.208333333332, 23762.211805555555, 23762.215277777777, 23762.21875, 23762.222222222223, 23762.225694444445, 23762.229166666668, 23762.23263888889, 23762.23611111111, 23762.239583333332, 23762.243055555555, 23762.246527777777, 23762.25, 23762.253472222223, 23762.256944444445, 23762.260416666668, 23762.26388888889, 23762.26736111111, 23762.270833333332, 23762.274305555555, 23762.277777777777, 23762.28125, 23762.284722222223, 23762.288194444445, 23762.291666666668, 23762.29513888889, 23762.29861111111, 23762.302083333332, 23762.305555555555, 23762.309027777777, 23762.3125, 23762.315972222223, 23762.319444444445, 23762.322916666668, 23762.32638888889, 23762.32986111111, 23762.333333333332, 23762.336805555555, 23762.340277777777, 23762.34375, 23762.347222222223, 23762.350694444445, 23762.354166666668, 23762.35763888889, 23762.36111111111, 23762.364583333332, 23762.368055555555, 23762.371527777777, 23762.375, 23762.378472222223, 23762.381944444445, 23762.385416666668, 23762.38888888889, 23762.39236111111, 23762.395833333332, 23762.399305555555, 23762.402777777777, 23762.40625, 23762.409722222223, 23762.413194444445, 23762.416666666668, 23762.42013888889, 23762.42361111111, 23762.427083333332, 23762.430555555555, 23762.434027777777, 23762.4375, 23762.440972222223, 23762.444444444445, 23762.447916666668, 23762.45138888889, 23762.45486111111, 23762.458333333332, 23762.461805555555, 23762.465277777777, 23762.46875, 23762.472222222223, 23762.475694444445, 23762.479166666668, 23762.48263888889, 23762.48611111111, 23762.489583333332, 23762.493055555555, 23762.496527777777, 23762.5, 23762.503472222223, 23762.506944444445, 23762.510416666668, 23762.51388888889, 23762.51736111111, 23762.520833333332, 23762.524305555555, 23762.527777777777, 23762.53125, 23762.534722222223, 23762.538194444445, 23762.541666666668, 23762.54513888889, 23762.54861111111, 23762.552083333332, 23762.555555555555, 23762.559027777777, 23762.5625, 23762.565972222223, 23762.569444444445, 23762.572916666668, 23762.57638888889, 23762.57986111111, 23762.583333333332, 23762.586805555555, 23762.590277777777, 23762.59375, 23762.597222222223, 23762.600694444445, 23762.604166666668, 23762.60763888889, 23762.61111111111, 23762.614583333332, 23762.618055555555, 23762.621527777777, 23762.625, 23762.628472222223, 23762.631944444445, 23762.635416666668, 23762.63888888889, 23762.64236111111, 23762.645833333332, 23762.649305555555, 23762.652777777777, 23762.65625, 23762.659722222223, 23762.663194444445, 23762.666666666668, 23762.67013888889, 23762.67361111111, 23762.677083333332, 23762.680555555555, 23762.684027777777, 23762.6875, 23762.690972222223, 23762.694444444445, 23762.697916666668, 23762.70138888889, 23762.70486111111, 23762.708333333332, 23762.711805555555, 23762.715277777777, 23762.71875, 23762.722222222223, 23762.725694444445, 23762.729166666668, 23762.73263888889, 23762.73611111111, 23762.739583333332, 23762.743055555555, 23762.746527777777, 23762.75, 23762.753472222223, 23762.756944444445, 23762.760416666668, 23762.76388888889, 23762.76736111111, 23762.770833333332, 23762.774305555555, 23762.777777777777, 23762.78125, 23762.784722222223, 23762.788194444445, 23762.791666666668, 23762.79513888889, 23762.79861111111, 23762.802083333332, 23762.805555555555, 23762.809027777777, 23762.8125, 23762.815972222223, 23762.819444444445, 23762.822916666668, 23762.82638888889, 23762.82986111111, 23762.833333333332, 23762.836805555555, 23762.840277777777, 23762.84375, 23762.847222222223, 23762.850694444445, 23762.854166666668, 23762.85763888889, 23762.86111111111, 23762.864583333332, 23762.868055555555, 23762.871527777777, 23762.875, 23762.878472222223, 23762.881944444445, 23762.885416666668, 23762.88888888889, 23762.89236111111, 23762.895833333332, 23762.899305555555, 23762.902777777777, 23762.90625, 23762.909722222223, 23762.913194444445, 23762.916666666668, 23762.92013888889, 23762.92361111111, 23762.927083333332, 23762.930555555555, 23762.934027777777, 23762.9375, 23762.940972222223, 23762.944444444445, 23762.947916666668, 23762.95138888889, 23762.95486111111, 23762.958333333332, 23762.961805555555, 23762.965277777777, 23762.96875, 23762.972222222223, 23762.975694444445, 23762.979166666668, 23762.98263888889, 23762.98611111111, 23762.989583333332, 23762.993055555555, 23762.996527777777, 23763.0, 23763.003472222223, 23763.006944444445, 23763.010416666668, 23763.01388888889, 23763.01736111111, 23763.020833333332, 23763.024305555555, 23763.027777777777, 23763.03125, 23763.034722222223, 23763.038194444445, 23763.041666666668, 23763.04513888889, 23763.04861111111, 23763.052083333332, 23763.055555555555, 23763.059027777777, 23763.0625, 23763.065972222223, 23763.069444444445, 23763.072916666668, 23763.07638888889, 23763.07986111111, 23763.083333333332, 23763.086805555555, 23763.090277777777, 23763.09375, 23763.097222222223, 23763.100694444445, 23763.104166666668, 23763.10763888889, 23763.11111111111, 23763.114583333332, 23763.118055555555, 23763.121527777777, 23763.125, 23763.128472222223, 23763.131944444445, 23763.135416666668, 23763.13888888889, 23763.14236111111, 23763.145833333332, 23763.149305555555, 23763.152777777777, 23763.15625, 23763.159722222223, 23763.163194444445, 23763.166666666668, 23763.17013888889, 23763.17361111111, 23763.177083333332, 23763.180555555555, 23763.184027777777, 23763.1875, 23763.190972222223, 23763.194444444445, 23763.197916666668, 23763.20138888889, 23763.20486111111, 23763.208333333332, 23763.211805555555, 23763.215277777777, 23763.21875, 23763.222222222223, 23763.225694444445, 23763.229166666668, 23763.23263888889, 23763.23611111111, 23763.239583333332, 23763.243055555555, 23763.246527777777, 23763.25, 23763.253472222223, 23763.256944444445, 23763.260416666668, 23763.26388888889, 23763.26736111111, 23763.270833333332, 23763.274305555555, 23763.277777777777, 23763.28125, 23763.284722222223, 23763.288194444445, 23763.291666666668, 23763.29513888889, 23763.29861111111, 23763.302083333332, 23763.305555555555, 23763.309027777777, 23763.3125, 23763.315972222223, 23763.319444444445, 23763.322916666668, 23763.32638888889, 23763.32986111111, 23763.333333333332, 23763.336805555555, 23763.340277777777, 23763.34375, 23763.347222222223, 23763.350694444445, 23763.354166666668, 23763.35763888889, 23763.36111111111, 23763.364583333332, 23763.368055555555, 23763.371527777777, 23763.375, 23763.378472222223, 23763.381944444445, 23763.385416666668, 23763.38888888889, 23763.39236111111, 23763.395833333332, 23763.399305555555, 23763.402777777777, 23763.40625, 23763.409722222223, 23763.413194444445, 23763.416666666668, 23763.42013888889, 23763.42361111111, 23763.427083333332, 23763.430555555555, 23763.434027777777, 23763.4375, 23763.440972222223, 23763.444444444445, 23763.447916666668, 23763.45138888889, 23763.45486111111, 23763.458333333332, 23763.461805555555, 23763.465277777777, 23763.46875, 23763.472222222223, 23763.475694444445, 23763.479166666668, 23763.48263888889, 23763.48611111111, 23763.489583333332, 23763.493055555555, 23763.496527777777, 23763.5, 23763.503472222223, 23763.506944444445, 23763.510416666668, 23763.51388888889, 23763.51736111111, 23763.520833333332, 23763.524305555555, 23763.527777777777, 23763.53125, 23763.534722222223, 23763.538194444445, 23763.541666666668, 23763.54513888889, 23763.54861111111, 23763.552083333332, 23763.555555555555, 23763.559027777777, 23763.5625, 23763.565972222223, 23763.569444444445, 23763.572916666668, 23763.57638888889, 23763.57986111111, 23763.583333333332, 23763.586805555555, 23763.590277777777, 23763.59375, 23763.597222222223, 23763.600694444445, 23763.604166666668, 23763.60763888889, 23763.61111111111, 23763.614583333332, 23763.618055555555, 23763.621527777777, 23763.625, 23763.628472222223, 23763.631944444445, 23763.635416666668, 23763.63888888889, 23763.64236111111, 23763.645833333332, 23763.649305555555, 23763.652777777777, 23763.65625, 23763.659722222223, 23763.663194444445, 23763.666666666668, 23763.67013888889, 23763.67361111111, 23763.677083333332, 23763.680555555555, 23763.684027777777, 23763.6875, 23763.690972222223, 23763.694444444445, 23763.697916666668, 23763.70138888889, 23763.70486111111, 23763.708333333332, 23763.711805555555, 23763.715277777777, 23763.71875, 23763.722222222223, 23763.725694444445, 23763.729166666668, 23763.73263888889, 23763.73611111111, 23763.739583333332, 23763.743055555555, 23763.746527777777, 23763.75, 23763.753472222223, 23763.756944444445, 23763.760416666668, 23763.76388888889, 23763.76736111111, 23763.770833333332, 23763.774305555555, 23763.777777777777, 23763.78125, 23763.784722222223, 23763.788194444445, 23763.791666666668, 23763.79513888889, 23763.79861111111, 23763.802083333332, 23763.805555555555, 23763.809027777777, 23763.8125, 23763.815972222223, 23763.819444444445, 23763.822916666668, 23763.82638888889, 23763.82986111111, 23763.833333333332, 23763.836805555555, 23763.840277777777, 23763.84375, 23763.847222222223, 23763.850694444445, 23763.854166666668, 23763.85763888889, 23763.86111111111, 23763.864583333332, 23763.868055555555, 23763.871527777777, 23763.875, 23763.878472222223, 23763.881944444445, 23763.885416666668, 23763.88888888889, 23763.89236111111, 23763.895833333332, 23763.899305555555, 23763.902777777777, 23763.90625, 23763.909722222223, 23763.913194444445, 23763.916666666668, 23763.92013888889, 23763.92361111111, 23763.927083333332, 23763.930555555555, 23763.934027777777, 23763.9375, 23763.940972222223, 23763.944444444445, 23763.947916666668, 23763.95138888889, 23763.95486111111, 23763.958333333332, 23763.961805555555, 23763.965277777777, 23763.96875, 23763.972222222223, 23763.975694444445, 23763.979166666668, 23763.98263888889, 23763.98611111111, 23763.989583333332, 23763.993055555555, 23763.996527777777, 23764.0, 23764.003472222223, 23764.006944444445, 23764.010416666668, 23764.01388888889, 23764.01736111111, 23764.020833333332, 23764.024305555555, 23764.027777777777, 23764.03125, 23764.034722222223, 23764.038194444445, 23764.041666666668, 23764.04513888889, 23764.04861111111, 23764.052083333332, 23764.055555555555, 23764.059027777777, 23764.0625, 23764.065972222223, 23764.069444444445, 23764.072916666668, 23764.07638888889, 23764.07986111111, 23764.083333333332, 23764.086805555555, 23764.090277777777, 23764.09375, 23764.097222222223, 23764.100694444445, 23764.104166666668, 23764.10763888889, 23764.11111111111, 23764.114583333332, 23764.118055555555, 23764.121527777777, 23764.125, 23764.128472222223, 23764.131944444445, 23764.135416666668, 23764.13888888889, 23764.14236111111, 23764.145833333332, 23764.149305555555, 23764.152777777777, 23764.15625, 23764.159722222223, 23764.163194444445, 23764.166666666668, 23764.17013888889, 23764.17361111111, 23764.177083333332, 23764.180555555555, 23764.184027777777, 23764.1875, 23764.190972222223, 23764.194444444445, 23764.197916666668, 23764.20138888889, 23764.20486111111, 23764.208333333332, 23764.211805555555, 23764.215277777777, 23764.21875, 23764.222222222223, 23764.225694444445, 23764.229166666668, 23764.23263888889, 23764.23611111111, 23764.239583333332, 23764.243055555555, 23764.246527777777, 23764.25, 23764.253472222223, 23764.256944444445, 23764.260416666668, 23764.26388888889, 23764.26736111111, 23764.270833333332, 23764.274305555555, 23764.277777777777, 23764.28125, 23764.284722222223, 23764.288194444445, 23764.291666666668, 23764.29513888889, 23764.29861111111, 23764.302083333332, 23764.305555555555, 23764.309027777777, 23764.3125, 23764.315972222223, 23764.319444444445, 23764.322916666668, 23764.32638888889, 23764.32986111111, 23764.333333333332, 23764.336805555555, 23764.340277777777, 23764.34375, 23764.347222222223, 23764.350694444445, 23764.354166666668, 23764.35763888889, 23764.36111111111, 23764.364583333332, 23764.368055555555, 23764.371527777777, 23764.375, 23764.378472222223, 23764.381944444445, 23764.385416666668, 23764.38888888889, 23764.39236111111, 23764.395833333332, 23764.399305555555, 23764.402777777777, 23764.40625, 23764.409722222223, 23764.413194444445, 23764.416666666668, 23764.42013888889, 23764.42361111111, 23764.427083333332, 23764.430555555555, 23764.434027777777, 23764.4375, 23764.440972222223, 23764.444444444445, 23764.447916666668, 23764.45138888889, 23764.45486111111, 23764.458333333332, 23764.461805555555, 23764.465277777777, 23764.46875, 23764.472222222223, 23764.475694444445, 23764.479166666668, 23764.48263888889, 23764.48611111111, 23764.489583333332, 23764.493055555555, 23764.496527777777, 23764.5, 23764.503472222223, 23764.506944444445, 23764.510416666668, 23764.51388888889, 23764.51736111111, 23764.520833333332, 23764.524305555555, 23764.527777777777, 23764.53125, 23764.534722222223, 23764.538194444445, 23764.541666666668, 23764.54513888889, 23764.54861111111, 23764.552083333332, 23764.555555555555, 23764.559027777777, 23764.5625, 23764.565972222223, 23764.569444444445, 23764.572916666668, 23764.57638888889, 23764.57986111111, 23764.583333333332, 23764.586805555555, 23764.590277777777, 23764.59375, 23764.597222222223, 23764.600694444445, 23764.604166666668, 23764.60763888889, 23764.61111111111, 23764.614583333332, 23764.618055555555, 23764.621527777777, 23764.625, 23764.628472222223, 23764.631944444445, 23764.635416666668, 23764.63888888889, 23764.64236111111, 23764.645833333332, 23764.649305555555, 23764.652777777777, 23764.65625, 23764.659722222223, 23764.663194444445, 23764.666666666668, 23764.67013888889, 23764.67361111111, 23764.677083333332, 23764.680555555555, 23764.684027777777, 23764.6875, 23764.690972222223, 23764.694444444445, 23764.697916666668, 23764.70138888889, 23764.70486111111, 23764.708333333332, 23764.711805555555, 23764.715277777777, 23764.71875, 23764.722222222223, 23764.725694444445, 23764.729166666668, 23764.73263888889, 23764.73611111111, 23764.739583333332, 23764.743055555555, 23764.746527777777, 23764.75, 23764.753472222223, 23764.756944444445, 23764.760416666668, 23764.76388888889, 23764.76736111111, 23764.770833333332, 23764.774305555555, 23764.777777777777, 23764.78125, 23764.784722222223, 23764.788194444445, 23764.791666666668, 23764.79513888889, 23764.79861111111, 23764.802083333332, 23764.805555555555, 23764.809027777777, 23764.8125, 23764.815972222223, 23764.819444444445, 23764.822916666668, 23764.82638888889, 23764.82986111111, 23764.833333333332, 23764.836805555555, 23764.840277777777, 23764.84375, 23764.847222222223, 23764.850694444445, 23764.854166666668, 23764.85763888889, 23764.86111111111, 23764.864583333332, 23764.868055555555, 23764.871527777777, 23764.875, 23764.878472222223, 23764.881944444445, 23764.885416666668, 23764.88888888889, 23764.89236111111, 23764.895833333332, 23764.899305555555, 23764.902777777777, 23764.90625, 23764.909722222223, 23764.913194444445, 23764.916666666668, 23764.92013888889, 23764.92361111111, 23764.927083333332, 23764.930555555555, 23764.934027777777, 23764.9375, 23764.940972222223, 23764.944444444445, 23764.947916666668, 23764.95138888889, 23764.95486111111, 23764.958333333332, 23764.961805555555, 23764.965277777777, 23764.96875, 23764.972222222223, 23764.975694444445, 23764.979166666668, 23764.98263888889, 23764.98611111111, 23764.989583333332, 23764.993055555555, 23764.996527777777, 23765.0, 23765.003472222223, 23765.006944444445, 23765.010416666668, 23765.01388888889, 23765.01736111111, 23765.020833333332, 23765.024305555555, 23765.027777777777, 23765.03125, 23765.034722222223, 23765.038194444445, 23765.041666666668, 23765.04513888889, 23765.04861111111, 23765.052083333332, 23765.055555555555, 23765.059027777777, 23765.0625, 23765.065972222223, 23765.069444444445, 23765.072916666668, 23765.07638888889, 23765.07986111111, 23765.083333333332, 23765.086805555555, 23765.090277777777, 23765.09375, 23765.097222222223, 23765.100694444445, 23765.104166666668, 23765.10763888889, 23765.11111111111, 23765.114583333332, 23765.118055555555, 23765.121527777777, 23765.125, 23765.128472222223, 23765.131944444445, 23765.135416666668, 23765.13888888889, 23765.14236111111, 23765.145833333332, 23765.149305555555, 23765.152777777777, 23765.15625, 23765.159722222223, 23765.163194444445, 23765.166666666668, 23765.17013888889, 23765.17361111111, 23765.177083333332, 23765.180555555555, 23765.184027777777, 23765.1875, 23765.190972222223, 23765.194444444445, 23765.197916666668, 23765.20138888889, 23765.20486111111, 23765.208333333332, 23765.211805555555, 23765.215277777777, 23765.21875, 23765.222222222223, 23765.225694444445, 23765.229166666668, 23765.23263888889, 23765.23611111111, 23765.239583333332, 23765.243055555555, 23765.246527777777, 23765.25, 23765.253472222223, 23765.256944444445, 23765.260416666668, 23765.26388888889, 23765.26736111111, 23765.270833333332, 23765.274305555555, 23765.277777777777, 23765.28125, 23765.284722222223, 23765.288194444445, 23765.291666666668, 23765.29513888889, 23765.29861111111, 23765.302083333332, 23765.305555555555, 23765.309027777777, 23765.3125, 23765.315972222223, 23765.319444444445, 23765.322916666668, 23765.32638888889, 23765.32986111111, 23765.333333333332, 23765.336805555555, 23765.340277777777, 23765.34375, 23765.347222222223, 23765.350694444445, 23765.354166666668, 23765.35763888889, 23765.36111111111, 23765.364583333332, 23765.368055555555, 23765.371527777777, 23765.375, 23765.378472222223, 23765.381944444445, 23765.385416666668, 23765.38888888889, 23765.39236111111, 23765.395833333332, 23765.399305555555, 23765.402777777777, 23765.40625, 23765.409722222223, 23765.413194444445, 23765.416666666668, 23765.42013888889, 23765.42361111111, 23765.427083333332, 23765.430555555555, 23765.434027777777, 23765.4375, 23765.440972222223, 23765.444444444445, 23765.447916666668, 23765.45138888889, 23765.45486111111, 23765.458333333332, 23765.461805555555, 23765.465277777777, 23765.46875, 23765.472222222223, 23765.475694444445, 23765.479166666668, 23765.48263888889, 23765.48611111111, 23765.489583333332, 23765.493055555555, 23765.496527777777, 23765.5, 23765.503472222223, 23765.506944444445, 23765.510416666668, 23765.51388888889, 23765.51736111111, 23765.520833333332, 23765.524305555555, 23765.527777777777, 23765.53125, 23765.534722222223, 23765.538194444445, 23765.541666666668, 23765.54513888889, 23765.54861111111, 23765.552083333332, 23765.555555555555, 23765.559027777777, 23765.5625, 23765.565972222223, 23765.569444444445, 23765.572916666668, 23765.57638888889, 23765.57986111111, 23765.583333333332, 23765.586805555555, 23765.590277777777, 23765.59375, 23765.597222222223, 23765.600694444445, 23765.604166666668, 23765.60763888889, 23765.61111111111, 23765.614583333332, 23765.618055555555, 23765.621527777777, 23765.625, 23765.628472222223, 23765.631944444445, 23765.635416666668, 23765.63888888889, 23765.64236111111, 23765.645833333332, 23765.649305555555, 23765.652777777777, 23765.65625, 23765.659722222223, 23765.663194444445, 23765.666666666668, 23765.67013888889, 23765.67361111111, 23765.677083333332, 23765.680555555555, 23765.684027777777, 23765.6875, 23765.690972222223, 23765.694444444445, 23765.697916666668, 23765.70138888889, 23765.70486111111, 23765.708333333332, 23765.711805555555, 23765.715277777777, 23765.71875, 23765.722222222223, 23765.725694444445, 23765.729166666668, 23765.73263888889, 23765.73611111111, 23765.739583333332, 23765.743055555555, 23765.746527777777, 23765.75, 23765.753472222223, 23765.756944444445, 23765.760416666668, 23765.76388888889, 23765.76736111111, 23765.770833333332, 23765.774305555555, 23765.777777777777, 23765.78125, 23765.784722222223, 23765.788194444445, 23765.791666666668, 23765.79513888889, 23765.79861111111, 23765.802083333332, 23765.805555555555, 23765.809027777777, 23765.8125, 23765.815972222223, 23765.819444444445, 23765.822916666668, 23765.82638888889, 23765.82986111111, 23765.833333333332, 23765.836805555555, 23765.840277777777, 23765.84375, 23765.847222222223, 23765.850694444445, 23765.854166666668, 23765.85763888889, 23765.86111111111, 23765.864583333332, 23765.868055555555, 23765.871527777777, 23765.875, 23765.878472222223, 23765.881944444445, 23765.885416666668, 23765.88888888889, 23765.89236111111, 23765.895833333332, 23765.899305555555, 23765.902777777777, 23765.90625, 23765.909722222223, 23765.913194444445, 23765.916666666668, 23765.92013888889, 23765.92361111111, 23765.927083333332, 23765.930555555555, 23765.934027777777, 23765.9375, 23765.940972222223, 23765.944444444445, 23765.947916666668, 23765.95138888889, 23765.95486111111, 23765.958333333332, 23765.961805555555, 23765.965277777777, 23765.96875, 23765.972222222223, 23765.975694444445, 23765.979166666668, 23765.98263888889, 23765.98611111111, 23765.989583333332, 23765.993055555555, 23765.996527777777, 23766.0, 23766.003472222223, 23766.006944444445, 23766.010416666668, 23766.01388888889, 23766.01736111111, 23766.020833333332, 23766.024305555555, 23766.027777777777, 23766.03125, 23766.034722222223, 23766.038194444445, 23766.041666666668, 23766.04513888889, 23766.04861111111, 23766.052083333332, 23766.055555555555, 23766.059027777777, 23766.0625, 23766.065972222223, 23766.069444444445, 23766.072916666668, 23766.07638888889, 23766.07986111111, 23766.083333333332, 23766.086805555555, 23766.090277777777, 23766.09375, 23766.097222222223, 23766.100694444445, 23766.104166666668, 23766.10763888889, 23766.11111111111, 23766.114583333332, 23766.118055555555, 23766.121527777777, 23766.125, 23766.128472222223, 23766.131944444445, 23766.135416666668, 23766.13888888889, 23766.14236111111, 23766.145833333332, 23766.149305555555, 23766.152777777777, 23766.15625, 23766.159722222223, 23766.163194444445, 23766.166666666668, 23766.17013888889, 23766.17361111111, 23766.177083333332, 23766.180555555555, 23766.184027777777, 23766.1875, 23766.190972222223, 23766.194444444445, 23766.197916666668, 23766.20138888889, 23766.20486111111, 23766.208333333332, 23766.211805555555, 23766.215277777777, 23766.21875, 23766.222222222223, 23766.225694444445, 23766.229166666668, 23766.23263888889, 23766.23611111111, 23766.239583333332, 23766.243055555555, 23766.246527777777, 23766.25, 23766.253472222223, 23766.256944444445, 23766.260416666668, 23766.26388888889, 23766.26736111111, 23766.270833333332, 23766.274305555555, 23766.277777777777, 23766.28125, 23766.284722222223, 23766.288194444445, 23766.291666666668, 23766.29513888889, 23766.29861111111, 23766.302083333332, 23766.305555555555, 23766.309027777777, 23766.3125, 23766.315972222223, 23766.319444444445, 23766.322916666668, 23766.32638888889, 23766.32986111111, 23766.333333333332, 23766.336805555555, 23766.340277777777, 23766.34375, 23766.347222222223, 23766.350694444445, 23766.354166666668, 23766.35763888889, 23766.36111111111, 23766.364583333332, 23766.368055555555, 23766.371527777777, 23766.375, 23766.378472222223, 23766.381944444445, 23766.385416666668, 23766.38888888889, 23766.39236111111, 23766.395833333332, 23766.399305555555, 23766.402777777777, 23766.40625, 23766.409722222223, 23766.413194444445, 23766.416666666668, 23766.42013888889, 23766.42361111111, 23766.427083333332, 23766.430555555555, 23766.434027777777, 23766.4375, 23766.440972222223, 23766.444444444445, 23766.447916666668, 23766.45138888889, 23766.45486111111, 23766.458333333332, 23766.461805555555, 23766.465277777777, 23766.46875, 23766.472222222223, 23766.475694444445, 23766.479166666668, 23766.48263888889, 23766.48611111111, 23766.489583333332, 23766.493055555555, 23766.496527777777, 23766.5, 23766.503472222223, 23766.506944444445, 23766.510416666668, 23766.51388888889, 23766.51736111111, 23766.520833333332, 23766.524305555555, 23766.527777777777, 23766.53125, 23766.534722222223, 23766.538194444445, 23766.541666666668, 23766.54513888889, 23766.54861111111, 23766.552083333332, 23766.555555555555, 23766.559027777777, 23766.5625, 23766.565972222223, 23766.569444444445, 23766.572916666668, 23766.57638888889, 23766.57986111111, 23766.583333333332, 23766.586805555555, 23766.590277777777, 23766.59375, 23766.597222222223, 23766.600694444445, 23766.604166666668, 23766.60763888889, 23766.61111111111, 23766.614583333332, 23766.618055555555, 23766.621527777777, 23766.625, 23766.628472222223, 23766.631944444445, 23766.635416666668, 23766.63888888889, 23766.64236111111, 23766.645833333332, 23766.649305555555, 23766.652777777777, 23766.65625, 23766.659722222223, 23766.663194444445, 23766.666666666668, 23766.67013888889, 23766.67361111111, 23766.677083333332, 23766.680555555555, 23766.684027777777, 23766.6875, 23766.690972222223, 23766.694444444445, 23766.697916666668, 23766.70138888889, 23766.70486111111, 23766.708333333332, 23766.711805555555, 23766.715277777777, 23766.71875, 23766.722222222223, 23766.725694444445, 23766.729166666668, 23766.73263888889, 23766.73611111111, 23766.739583333332, 23766.743055555555, 23766.746527777777, 23766.75, 23766.753472222223, 23766.756944444445, 23766.760416666668, 23766.76388888889, 23766.76736111111, 23766.770833333332, 23766.774305555555, 23766.777777777777, 23766.78125, 23766.784722222223, 23766.788194444445, 23766.791666666668, 23766.79513888889, 23766.79861111111, 23766.802083333332, 23766.805555555555, 23766.809027777777, 23766.8125, 23766.815972222223, 23766.819444444445, 23766.822916666668, 23766.82638888889, 23766.82986111111, 23766.833333333332, 23766.836805555555, 23766.840277777777, 23766.84375, 23766.847222222223, 23766.850694444445, 23766.854166666668, 23766.85763888889, 23766.86111111111, 23766.864583333332, 23766.868055555555, 23766.871527777777, 23766.875, 23766.878472222223, 23766.881944444445, 23766.885416666668, 23766.88888888889, 23766.89236111111, 23766.895833333332, 23766.899305555555, 23766.902777777777, 23766.90625, 23766.909722222223, 23766.913194444445, 23766.916666666668, 23766.92013888889, 23766.92361111111, 23766.927083333332, 23766.930555555555, 23766.934027777777, 23766.9375, 23766.940972222223, 23766.944444444445, 23766.947916666668, 23766.95138888889, 23766.95486111111, 23766.958333333332, 23766.961805555555, 23766.965277777777, 23766.96875, 23766.972222222223, 23766.975694444445, 23766.979166666668, 23766.98263888889, 23766.98611111111, 23766.989583333332, 23766.993055555555, 23766.996527777777, 23767.0, 23767.003472222223, 23767.006944444445, 23767.010416666668, 23767.01388888889, 23767.01736111111, 23767.020833333332, 23767.024305555555, 23767.027777777777, 23767.03125, 23767.034722222223, 23767.038194444445, 23767.041666666668, 23767.04513888889, 23767.04861111111, 23767.052083333332, 23767.055555555555, 23767.059027777777, 23767.0625, 23767.065972222223, 23767.069444444445, 23767.072916666668, 23767.07638888889, 23767.07986111111, 23767.083333333332, 23767.086805555555, 23767.090277777777, 23767.09375, 23767.097222222223, 23767.100694444445, 23767.104166666668, 23767.10763888889, 23767.11111111111, 23767.114583333332, 23767.118055555555, 23767.121527777777, 23767.125, 23767.128472222223, 23767.131944444445, 23767.135416666668, 23767.13888888889, 23767.14236111111, 23767.145833333332, 23767.149305555555, 23767.152777777777, 23767.15625, 23767.159722222223, 23767.163194444445, 23767.166666666668, 23767.17013888889, 23767.17361111111, 23767.177083333332, 23767.180555555555, 23767.184027777777, 23767.1875, 23767.190972222223, 23767.194444444445, 23767.197916666668, 23767.20138888889, 23767.20486111111, 23767.208333333332, 23767.211805555555, 23767.215277777777, 23767.21875, 23767.222222222223, 23767.225694444445, 23767.229166666668, 23767.23263888889, 23767.23611111111, 23767.239583333332, 23767.243055555555, 23767.246527777777, 23767.25, 23767.253472222223, 23767.256944444445, 23767.260416666668, 23767.26388888889, 23767.26736111111, 23767.270833333332, 23767.274305555555, 23767.277777777777, 23767.28125, 23767.284722222223, 23767.288194444445, 23767.291666666668, 23767.29513888889, 23767.29861111111, 23767.302083333332, 23767.305555555555, 23767.309027777777, 23767.3125, 23767.315972222223, 23767.319444444445, 23767.322916666668, 23767.32638888889, 23767.32986111111, 23767.333333333332, 23767.336805555555, 23767.340277777777, 23767.34375, 23767.347222222223, 23767.350694444445, 23767.354166666668, 23767.35763888889, 23767.36111111111, 23767.364583333332, 23767.368055555555, 23767.371527777777, 23767.375, 23767.378472222223, 23767.381944444445, 23767.385416666668, 23767.38888888889, 23767.39236111111, 23767.395833333332, 23767.399305555555, 23767.402777777777, 23767.40625, 23767.409722222223, 23767.413194444445, 23767.416666666668, 23767.42013888889, 23767.42361111111, 23767.427083333332, 23767.430555555555, 23767.434027777777, 23767.4375, 23767.440972222223, 23767.444444444445, 23767.447916666668, 23767.45138888889, 23767.45486111111, 23767.458333333332, 23767.461805555555, 23767.465277777777, 23767.46875, 23767.472222222223, 23767.475694444445, 23767.479166666668, 23767.48263888889, 23767.48611111111, 23767.489583333332, 23767.493055555555, 23767.496527777777, 23767.5, 23767.503472222223, 23767.506944444445, 23767.510416666668, 23767.51388888889, 23767.51736111111, 23767.520833333332, 23767.524305555555, 23767.527777777777, 23767.53125, 23767.534722222223, 23767.538194444445, 23767.541666666668, 23767.54513888889, 23767.54861111111, 23767.552083333332, 23767.555555555555, 23767.559027777777, 23767.5625, 23767.565972222223, 23767.569444444445, 23767.572916666668, 23767.57638888889, 23767.57986111111, 23767.583333333332, 23767.586805555555, 23767.590277777777, 23767.59375, 23767.597222222223, 23767.600694444445, 23767.604166666668, 23767.60763888889, 23767.61111111111, 23767.614583333332, 23767.618055555555, 23767.621527777777, 23767.625, 23767.628472222223, 23767.631944444445, 23767.635416666668, 23767.63888888889, 23767.64236111111, 23767.645833333332, 23767.649305555555, 23767.652777777777, 23767.65625, 23767.659722222223, 23767.663194444445, 23767.666666666668, 23767.67013888889, 23767.67361111111, 23767.677083333332, 23767.680555555555, 23767.684027777777, 23767.6875, 23767.690972222223, 23767.694444444445, 23767.697916666668, 23767.70138888889, 23767.70486111111, 23767.708333333332, 23767.711805555555, 23767.715277777777, 23767.71875, 23767.722222222223, 23767.725694444445, 23767.729166666668, 23767.73263888889, 23767.73611111111, 23767.739583333332, 23767.743055555555, 23767.746527777777, 23767.75, 23767.753472222223, 23767.756944444445, 23767.760416666668, 23767.76388888889, 23767.76736111111, 23767.770833333332, 23767.774305555555, 23767.777777777777, 23767.78125, 23767.784722222223, 23767.788194444445, 23767.791666666668, 23767.79513888889, 23767.79861111111, 23767.802083333332, 23767.805555555555, 23767.809027777777, 23767.8125, 23767.815972222223, 23767.819444444445, 23767.822916666668, 23767.82638888889, 23767.82986111111, 23767.833333333332, 23767.836805555555, 23767.840277777777, 23767.84375, 23767.847222222223, 23767.850694444445, 23767.854166666668, 23767.85763888889, 23767.86111111111, 23767.864583333332, 23767.868055555555, 23767.871527777777, 23767.875, 23767.878472222223, 23767.881944444445, 23767.885416666668, 23767.88888888889, 23767.89236111111, 23767.895833333332, 23767.899305555555, 23767.902777777777, 23767.90625, 23767.909722222223, 23767.913194444445, 23767.916666666668, 23767.92013888889, 23767.92361111111, 23767.927083333332, 23767.930555555555, 23767.934027777777, 23767.9375, 23767.940972222223, 23767.944444444445, 23767.947916666668, 23767.95138888889, 23767.95486111111, 23767.958333333332, 23767.961805555555, 23767.965277777777, 23767.96875, 23767.972222222223, 23767.975694444445, 23767.979166666668, 23767.98263888889, 23767.98611111111, 23767.989583333332, 23767.993055555555, 23767.996527777777, 23768.0, 23768.003472222223, 23768.006944444445, 23768.010416666668, 23768.01388888889, 23768.01736111111, 23768.020833333332, 23768.024305555555, 23768.027777777777, 23768.03125, 23768.034722222223, 23768.038194444445, 23768.041666666668, 23768.04513888889, 23768.04861111111, 23768.052083333332, 23768.055555555555, 23768.059027777777, 23768.0625, 23768.065972222223, 23768.069444444445, 23768.072916666668, 23768.07638888889, 23768.07986111111, 23768.083333333332, 23768.086805555555, 23768.090277777777, 23768.09375, 23768.097222222223, 23768.100694444445, 23768.104166666668, 23768.10763888889, 23768.11111111111, 23768.114583333332, 23768.118055555555, 23768.121527777777, 23768.125, 23768.128472222223, 23768.131944444445, 23768.135416666668, 23768.13888888889, 23768.14236111111, 23768.145833333332, 23768.149305555555, 23768.152777777777, 23768.15625, 23768.159722222223, 23768.163194444445, 23768.166666666668, 23768.17013888889, 23768.17361111111, 23768.177083333332, 23768.180555555555, 23768.184027777777, 23768.1875, 23768.190972222223, 23768.194444444445, 23768.197916666668, 23768.20138888889, 23768.20486111111, 23768.208333333332, 23768.211805555555, 23768.215277777777, 23768.21875, 23768.222222222223, 23768.225694444445, 23768.229166666668, 23768.23263888889, 23768.23611111111, 23768.239583333332, 23768.243055555555, 23768.246527777777, 23768.25, 23768.253472222223, 23768.256944444445, 23768.260416666668, 23768.26388888889}
LATITUDE =-31.9966
LONGITUDE =115.4157166667
NOMINAL_DEPTH =43.0
TEMP =
  {19.868317, 19.868008, 19.868235, 19.869808, 19.867914, 19.86762, 19.870531, 19.868395, 19.868607, 19.871466, 19.871145, 19.868755, 19.870562, 19.872295, 19.872585, 19.872126, 19.873642, 19.872622, 19.880365, 19.87585, 19.875381, 19.876574, 19.878492, 19.879908, 19.880716, 19.880154, 19.882643, 19.88546, 19.883993, 19.885412, 19.88614, 19.887587, 19.888918, 19.889935, 19.891272, 19.892727, 19.89381, 19.89495, 19.894243, 19.897568, 19.899761, 19.90199, 19.902699, 19.905016, 19.9061, 19.908468, 19.90717, 19.910002, 19.910013, 19.911112, 19.913214, 19.910452, 19.91594, 19.915295, 19.915232, 19.914824, 19.920292, 19.91897, 19.917953, 19.919945, 19.919672, 19.921406, 19.923178, 19.925259, 19.926039, 19.926756, 19.927431, 19.928686, 19.929832, 19.931093, 19.931976, 19.93341, 19.933546, 19.933706, 19.933943, 19.93544, 19.936138, 19.937346, 19.939474, 19.940239, 19.9422, 19.944262, 19.947556, 19.951496, 19.954792, 19.952747, 19.953918, 19.961496, 19.958923, 19.962276, 19.964369, 19.971048, 19.983938, 19.974958, 19.97329, 19.975233, 19.973682, 19.971233, 19.969297, 19.966316, 19.967281, 19.964714, 19.964327, 19.9582, 19.956894, 19.955666, 19.955862, 19.955923, 19.95599, 19.953619, 19.955954, 19.950495, 19.951384, 19.948042, 19.945892, 19.943708, 19.944302, 19.945562, 19.949993, 19.948816, 19.952255, 19.952887, 19.955065, 19.95947, 19.960783, 19.96176, 19.960447, 19.963171, 19.962452, 19.964659, 19.965721, 19.969818, 19.977402, 19.976461, 19.981127, 19.984285, 19.98631, 19.99048, 19.989468, 19.99142, 19.995104, 19.999868, 20.0139, 20.017385, 20.01493, 20.015663, 20.02564, 20.024979, 20.024508, 20.028236, 20.032413, 20.03204, 20.03536, 20.032728, 20.035086, 20.036978, 20.03991, 20.037195, 20.037909, 20.03855, 20.035086, 20.038897, 20.03628, 20.03916, 20.036715, 20.037779, 20.035717, 20.033783, 20.033333, 20.035173, 20.035128, 20.037775, 20.036388, 20.035702, 20.035183, 20.036673, 20.038364, 20.041115, 20.039362, 20.042034, 20.043715, 20.044724, 20.045183, 20.0466, 20.04778, 20.046326, 20.044832, 20.041155, 20.042929, 20.04218, 20.043787, 20.046305, 20.048792, 20.049429, 20.051352, 20.050209, 20.049221, 20.047567, 20.04828, 20.046331, 20.047861, 20.044376, 20.0463, 20.043224, 20.045395, 20.043566, 20.04099, 20.045359, 20.044724, 20.041466, 20.041864, 20.039062, 20.041409, 20.04188, 20.042593, 20.041016, 20.040438, 20.04399, 20.040127, 20.039885, 20.038824, 20.040033, 20.04094, 20.039326, 20.038757, 20.040846, 20.03659, 20.035654, 20.03478, 20.033602, 20.036192, 20.0331, 20.030376, 20.026457, 20.023954, 20.02444, 20.02444, 20.024565, 20.023129, 20.022694, 20.02244, 20.021898, 20.022135, 20.022348, 20.027046, 20.02506, 20.023273, 20.022549, 20.021402, 20.022709, 20.022306, 20.024084, 20.022736, 20.022425, 20.02227, 20.022648, 20.021065, 20.02256, 20.021872, 20.023035, 20.020922, 20.022709, 20.020306, 20.023117, 20.02212, 20.021872, 20.023216, 20.020493, 20.019976, 20.021261, 20.020203, 20.020332, 20.020502, 20.020182, 20.020327, 20.019102, 20.017908, 20.01922, 20.021536, 20.03128, 20.022947, 20.020777, 20.022875, 20.021019, 20.021923, 20.019794, 20.024141, 20.019701, 20.018703, 20.017872, 20.01751, 20.016998, 20.016802, 20.016672, 20.022053, 20.029129, 20.020472, 20.018978, 20.020704, 20.018135, 20.01797, 20.017763, 20.018265, 20.018208, 20.019323, 20.017706, 20.017654, 20.017664, 20.017979, 20.018063, 20.017199, 20.017235, 20.017323, 20.017174, 20.017736, 20.016212, 20.016518, 20.015778, 20.016155, 20.017065, 20.01711, 20.017767, 20.01845, 20.018677, 20.018894, 20.019133, 20.020704, 20.022135, 20.022793, 20.023685, 20.025024, 20.02642, 20.025108, 20.02682, 20.025843, 20.026545, 20.027775, 20.02883, 20.028793, 20.02928, 20.030128, 20.033901, 20.031202, 20.031958, 20.032686, 20.0337, 20.035189, 20.034605, 20.035505, 20.035732, 20.036192, 20.041176, 20.035355, 20.03822, 20.037918, 20.03945, 20.0398, 20.041786, 20.041864, 20.042402, 20.04311, 20.043037, 20.044191, 20.045395, 20.04641, 20.051756, 20.048819, 20.049238, 20.050365, 20.051647, 20.05159, 20.053467, 20.052113, 20.0519, 20.052412, 20.052874, 20.054708, 20.055473, 20.055883, 20.057041, 20.055065, 20.055593, 20.056223, 20.05566, 20.055836, 20.055561, 20.056679, 20.056498, 20.056488, 20.058023, 20.05809, 20.057894, 20.057129, 20.056803, 20.056684, 20.0477, 20.043037, 20.038782, 20.03704, 20.035355, 20.027336, 20.02456, 20.014336, 20.017887, 20.039656, 20.010738, 20.007229, 20.000004, 19.99631, 19.9928, 19.987518, 19.9817, 19.968218, 19.960773, 19.953102, 19.940042, 19.937454, 19.92056, 19.910173, 19.90495, 19.903969, 19.891342, 19.882084, 19.881817, 19.878998, 19.880604, 19.880903, 19.893335, 19.88354, 19.884335, 19.888546, 19.887865, 19.892437, 19.889288, 19.892065, 19.889763, 19.894869, 19.887657, 19.889835, 19.89041, 19.888025, 19.908062, 19.883472, 19.865469, 19.863478, 19.853825, 19.849106, 19.841888, 19.831789, 19.828236, 19.79983, 19.78199, 19.742378, 19.711899, 19.700817, 19.689083, 19.683306, 19.666956, 19.665943, 19.630322, 19.620562, 19.604408, 19.585663, 19.570845, 19.555534, 19.53281, 19.514883, 19.51145, 19.499855, 19.48543, 19.470875, 19.459969, 19.45165, 19.446115, 19.433596, 19.417175, 19.403263, 19.398018, 19.396223, 19.372879, 19.34765, 19.343964, 19.336958, 19.331217, 19.327192, 19.321178, 19.30644, 19.280575, 19.266525, 19.254286, 19.24237, 19.218807, 19.215895, 19.20032, 19.19226, 19.1795, 19.16734, 19.166904, 19.160196, 19.143015, 19.139555, 19.13753, 19.13263, 19.126572, 19.117712, 19.115166, 19.110256, 19.100176, 19.088385, 19.086231, 19.087091, 19.087719, 19.085577, 19.078543, 19.068993, 19.068287, 19.06408, 19.058565, 19.057056, 19.055206, 19.048119, 19.042885, 19.039455, 19.034254, 19.028284, 19.029001, 19.024862, 19.022486, 19.020693, 19.017643, 19.010597, 19.00745, 19.001244, 18.994062, 18.987804, 18.981115, 18.977331, 18.975605, 18.972284, 18.96919, 18.965662, 18.958897, 18.952755, 18.949411, 18.945246, 18.942299, 18.937088, 18.930748, 18.92813, 18.923643, 18.914953, 18.909027, 18.906069, 18.903261, 18.899231, 18.89737, 18.893282, 18.88563, 18.881319, 18.877289, 18.872437, 18.870148, 18.867525, 18.867031, 18.863771, 18.862038, 18.859905, 18.857355, 18.856785, 18.855244, 18.854208, 18.851746, 18.851532, 18.847248, 18.840715, 18.827679, 18.824516, 18.820683, 18.820265, 18.818935, 18.817268, 18.812786, 18.810804, 18.808954, 18.801262, 18.797766, 18.789234, 18.780077, 18.771088, 18.761908, 18.755856, 18.752249, 18.746946, 18.754078, 18.743406, 18.739988, 18.735796, 18.729734, 18.719275, 18.714325, 18.715868, 18.714325, 18.710806, 18.711391, 18.709152, 18.706179, 18.7046, 18.700165, 18.697075, 18.695543, 18.688553, 18.685686, 18.684374, 18.680637, 18.67287, 18.666868, 18.655195, 18.649317, 18.639898, 18.637524, 18.636465, 18.632029, 18.630146, 18.622814, 18.624397, 18.628487, 18.626152, 18.621681, 18.620266, 18.62046, 18.618963, 18.615892, 18.613445, 18.615469, 18.612728, 18.61433, 18.608276, 18.616152, 18.617245, 18.607769, 18.606167, 18.606537, 18.611975, 18.610836, 18.608877, 18.610235, 18.609737, 18.607204, 18.620623, 18.608038, 18.602205, 18.601091, 18.601076, 18.60024, 18.597937, 18.599264, 18.599865, 18.597301, 18.586693, 18.588697, 18.64288, 18.586693, 18.582722, 18.574938, 18.576315, 18.569456, 18.565094, 18.56394, 18.561623, 18.553509, 18.558273, 18.558765, 18.560081, 18.561293, 18.559843, 18.576956, 18.587528, 18.571781, 18.571007, 18.588148, 18.586678, 18.583652, 18.578, 18.578512, 18.584192, 18.59181, 18.568695, 18.59626, 18.59872, 18.598497, 18.59457, 18.58795, 18.631544, 18.59537, 18.594591, 18.597845, 18.593197, 18.594393, 18.605175, 18.592821, 18.587715, 18.595741, 18.590364, 18.582077, 18.573118, 18.579311, 18.568491, 18.571964, 18.572386, 18.5706, 18.567581, 18.563015, 18.555435, 18.55083, 18.546728, 18.540552, 18.535221, 18.54841, 18.534399, 18.537828, 18.544939, 18.546795, 18.540024, 18.534958, 18.532898, 18.529612, 18.527252, 18.527786, 18.527008, 18.530058, 18.528812, 18.536522, 18.541437, 18.541758, 18.528812, 18.52892, 18.526663, 18.52584, 18.528553, 18.527548, 18.534369, 18.53513, 18.537184, 18.540695, 18.546652, 18.532522, 18.52731, 18.535004, 18.523664, 18.537554, 18.518091, 18.512638, 18.508497, 18.508762, 18.50834, 18.510235, 18.515875, 18.51171, 18.511652, 18.511892, 18.511831, 18.513756, 18.511557, 18.514696, 18.511145, 18.510397, 18.510601, 18.510073, 18.510021, 18.510118, 18.509016, 18.511093, 18.507456, 18.502182, 18.496761, 18.491737, 18.488598, 18.486734, 18.48328, 18.478125, 18.47246, 18.468534, 18.471405, 18.465736, 18.46112, 18.459154, 18.454107, 18.443592, 18.43958, 18.432564, 18.42294, 18.420208, 18.407335, 18.396023, 18.388979, 18.3835, 18.381317, 18.378466, 18.379847, 18.374954, 18.367264, 18.35806, 18.355007, 18.348267, 18.349209, 18.351385, 18.350351, 18.345638, 18.347383, 18.343021, 18.340475, 18.336767, 18.33445, 18.33205, 18.331285, 18.326473, 18.324484, 18.317883, 18.314547, 18.316935, 18.31293, 18.315155, 18.313278, 18.312021, 18.31092, 18.310272, 18.314009, 18.310946, 18.312006, 18.311981, 18.308603, 18.306728, 18.305243, 18.302555, 18.299047, 18.296663, 18.295776, 18.297804, 18.29267, 18.289835, 18.288397, 18.288736, 18.294828, 18.30075, 18.296375, 18.29751, 18.30002, 18.300917, 18.296394, 18.29847, 18.296263, 18.304283, 18.298038, 18.29891, 18.299934, 18.29601, 18.29819, 18.295883, 18.295366, 18.294737, 18.29199, 18.29348, 18.292324, 18.30111, 18.298824, 18.298708, 18.304136, 18.304802, 18.30398, 18.319439, 18.307219, 18.307047, 18.303102, 18.30498, 18.30227, 18.300085, 18.303225, 18.309166, 18.322035, 18.318974, 18.318075, 18.3138, 18.319374, 18.314388, 18.311697, 18.309166, 18.303812, 18.30194, 18.323318, 18.310606, 18.307823, 18.309475, 18.305582, 18.299818, 18.288979, 18.288563, 18.28615, 18.281792, 18.280458, 18.278522, 18.27468, 18.273975, 18.276712, 18.281801, 18.271183, 18.27321, 18.271584, 18.27021, 18.27329, 18.275223, 18.280043, 18.279236, 18.281837, 18.27732, 18.28545, 18.285168, 18.307032, 18.292994, 18.284918, 18.286024, 18.283068, 18.280209, 18.28094, 18.285198, 18.280504, 18.286572, 18.293947, 18.287966, 18.303316, 18.28793, 18.294413, 18.29418, 18.308882, 18.309258, 18.301136, 18.31699, 18.303356, 18.303326, 18.30264, 18.311747, 18.304218, 18.314632, 18.32274, 18.321396, 18.32381, 18.324125, 18.322197, 18.323597, 18.32315, 18.343285, 18.320778, 18.314003, 18.31869, 18.31694, 18.330029, 18.32488, 18.324419, 18.330194, 18.325449, 18.323177, 18.319582, 18.31594, 18.309399, 18.30952, 18.323963, 18.298155, 18.29165, 18.28278, 18.275034, 18.276976, 18.27881, 18.279135, 18.282177, 18.272303, 18.268785, 18.265715, 18.261314, 18.25825, 18.254215, 18.254946, 18.245916, 18.245049, 18.23866, 18.242332, 18.23972, 18.226517, 18.224602, 18.220499, 18.218431, 18.217514, 18.215574, 18.211294, 18.211288, 18.213139, 18.214369, 18.220037, 18.214197, 18.21326, 18.210205, 18.209248, 18.209583, 18.208574, 18.2097, 18.207466, 18.211218, 18.210407, 18.213741, 18.21443, 18.212894, 18.215614, 18.234835, 18.213848, 18.214987, 18.213533, 18.22712, 18.217905, 18.222443, 18.216587, 18.21678, 18.225985, 18.221252, 18.215782, 18.220148, 18.228157, 18.215717, 18.233051, 18.222996, 18.22495, 18.216436, 18.217915, 18.210545, 18.200953, 18.201225, 18.200476, 18.199995, 18.202877, 18.19727, 18.19923, 18.204214, 18.200558, 18.197254, 18.200172, 18.194384, 18.193508, 18.189096, 18.200071, 18.193169, 18.190647, 18.19096, 18.192732, 18.197636, 18.197954, 18.197777, 18.210098, 18.19811, 18.19963, 18.195898, 18.196556, 18.208635, 18.201763, 18.20613, 18.199802, 18.205202, 18.20008, 18.201675, 18.2152, 18.199068, 18.206558, 18.207409, 18.20225, 18.199245, 18.200785, 18.204285, 18.204199, 18.212034, 18.207602, 18.211056, 18.209284, 18.205288, 18.207531, 18.209587, 18.209923, 18.214952, 18.218603, 18.220184, 18.217733, 18.218117, 18.217241, 18.217587, 18.215195, 18.215366, 18.21518, 18.216091, 18.218279, 18.214977, 18.21525, 18.216516, 18.216421, 18.21897, 18.215311, 18.217606, 18.216293, 18.216455, 18.216244, 18.21566, 18.21675, 18.216036, 18.217049, 18.216055, 18.21286, 18.212322, 18.2121, 18.211563, 18.206396, 18.205395, 18.202026, 18.20277, 18.201033, 18.201235, 18.19994, 18.200264, 18.197716, 18.191856, 18.19129, 18.189886, 18.190323, 18.18938, 18.1839, 18.184103, 18.183046, 18.181177, 18.180773, 18.180134, 18.179262, 18.176184, 18.175608, 18.170185, 18.17092, 18.16912, 18.169466, 18.171177, 18.168823, 18.168135, 18.167141, 18.167303, 18.167511, 18.16748, 18.167355, 18.165096, 18.165283, 18.162514, 18.163198, 18.164276, 18.165087, 18.164108, 18.163143, 18.163198, 18.165607, 18.164377, 18.164833, 18.164215, 18.164104, 18.164429, 18.165182, 18.164843, 18.165567, 18.165558, 18.166687, 18.167814, 18.169374, 18.170807, 18.171896, 18.171562, 18.172722, 18.172918, 18.173754, 18.174528, 18.17708, 18.177435, 18.178457, 18.180244, 18.182787, 18.183588, 18.183956, 18.185795, 18.18935, 18.188894, 18.193304, 18.193897, 18.195316, 18.201246, 18.20321, 18.206453, 18.20754, 18.209719, 18.214323, 18.21597, 18.214708, 18.214699, 18.21725, 18.21991, 18.219055, 18.220139, 18.224424, 18.222975, 18.223856, 18.227484, 18.22835, 18.230797, 18.230656, 18.232155, 18.232779, 18.236437, 18.236609, 18.241179, 18.245874, 18.24625, 18.246984, 18.256105, 18.252838, 18.255026, 18.254429, 18.259851, 18.257809, 18.264807, 18.272602, 18.265795, 18.271746, 18.269247, 18.27728, 18.276052, 18.282942, 18.283321, 18.288944, 18.29091, 18.297638, 18.301023, 18.304445, 18.329998, 18.347866, 18.340551, 18.33913, 18.363428, 18.444286, 18.409214, 18.556433, 18.570957, 18.584461, 18.606777, 18.663103, 18.662624, 18.660782, 18.697737, 18.706362, 18.718933, 18.779873, 18.728273, 18.745071, 18.738724, 18.750414, 18.712437, 18.680735, 18.684862, 18.665318, 18.665775, 18.634876, 18.65899, 18.611624, 18.672585, 18.62223, 18.655449, 18.624733, 18.67571, 18.638977, 18.658146, 18.67719, 18.649057, 18.691755, 18.71127, 18.708918, 18.708357, 18.709686, 18.711178, 18.714727, 18.711544, 18.725023, 18.723965, 18.724342, 18.72788, 18.736235, 18.73138, 18.740257, 18.737019, 18.74369, 18.741272, 18.737787, 18.74689, 18.694046, 18.74502, 18.74504, 18.686455, 18.737986, 18.675745, 18.75453, 18.747145, 18.725904, 18.743681, 18.745478, 18.773575, 18.787771, 18.785534, 18.781345, 18.782564, 18.782665, 18.780489, 18.779043, 18.779226, 18.78638, 18.78415, 18.783262, 18.783512, 18.774258, 18.771383, 18.761673, 18.748846, 18.751892, 18.727877, 18.727097, 18.71757, 18.717554, 18.702034, 18.69567, 18.683502, 18.681059, 18.670885, 18.66097, 18.65112, 18.647852, 18.642132, 18.635386, 18.63033, 18.629652, 18.62924, 18.626192, 18.62769, 18.62779, 18.629719, 18.627583, 18.626448, 18.626463, 18.625816, 18.625124, 18.62462, 18.626793, 18.627016, 18.62546, 18.622398, 18.623446, 18.622463, 18.622215, 18.62164, 18.619488, 18.62246, 18.622433, 18.619799, 18.6213, 18.621508, 18.622784, 18.624174, 18.62543, 18.62668, 18.627403, 18.63036, 18.631153, 18.63469, 18.634064, 18.634964, 18.640026, 18.637579, 18.639675, 18.644636, 18.645226, 18.648804, 18.64856, 18.650284, 18.657602, 18.656843, 18.656319, 18.659409, 18.660563, 18.666798, 18.67001, 18.67629, 18.673222, 18.67997, 18.685762, 18.684332, 18.68948, 18.690279, 18.692402, 18.693497, 18.702385, 18.707884, 18.714813, 18.71427, 18.715288, 18.722412, 18.724352, 18.73328, 18.730545, 18.733376, 18.73931, 18.740705, 18.741245, 18.74448, 18.742708, 18.752645, 18.74316, 18.74495, 18.74419, 18.748535, 18.749962, 18.754948, 18.76152, 18.76369, 18.763136, 18.7671, 18.77196, 18.772903, 18.774508, 18.777279, 18.777754, 18.784168, 18.785357, 18.791359, 18.796732, 18.7995, 18.80402, 18.808275, 18.813082, 18.81767, 18.823053, 18.83059, 18.836428, 18.842644, 18.845167, 18.845642, 18.848083, 18.854795, 18.855759, 18.857407, 18.862026, 18.864868, 18.867464, 18.870968, 18.874565, 18.881767, 18.882093, 18.886848, 18.894613, 18.900236, 18.908655, 18.914759, 18.916927, 18.920673, 18.92367, 18.932693, 18.9318, 18.935143, 18.93764, 18.947762, 18.950937, 18.954205, 18.957958, 18.95974, 18.96044, 18.966846, 18.968, 18.973434, 18.977222, 18.981197, 18.983862, 18.990961, 18.990313, 18.995268, 19.00205, 19.004288, 19.008364, 19.017994, 19.019793, 19.027584, 19.033466, 19.035791, 19.03919, 19.04249, 19.046917, 19.053383, 19.059225, 19.065071, 19.06798, 19.070505, 19.074223, 19.076635, 19.077335, 19.080608, 19.084837, 19.089136, 19.087362, 19.0893, 19.094894, 19.092598, 19.096565, 19.096382, 19.102335, 19.10267, 19.10508, 19.106302, 19.109667, 19.113283, 19.111954, 19.111048, 19.115314, 19.117073, 19.119226, 19.122623, 19.122828, 19.12419, 19.127094, 19.1296, 19.133877, 19.132986, 19.134676, 19.135626, 19.135555, 19.139597, 19.142212, 19.142082, 19.145823, 19.145302, 19.149343, 19.150269, 19.148024, 19.14833, 19.147516, 19.148914, 19.149317, 19.145828, 19.145357, 19.148167, 19.147379, 19.146591, 19.159117, 19.153719, 19.152914, 19.154772, 19.157024, 19.155994, 19.157715, 19.159372, 19.161184, 19.161716, 19.163006, 19.16668, 19.17141, 19.171383, 19.173025, 19.175402, 19.17768, 19.178312, 19.183954, 19.192871, 19.180412, 19.180176, 19.181221, 19.179604, 19.17974, 19.182106, 19.182648, 19.183842, 19.181768, 19.187016, 19.189974, 19.188044, 19.194729, 19.196583, 19.204493, 19.202951, 19.204575, 19.209044, 19.206749, 19.210594, 19.211634, 19.212904, 19.222588, 19.228952, 19.229618, 19.235477, 19.245798, 19.252806, 19.256018, 19.26057, 19.262707, 19.26381, 19.265839, 19.263123, 19.266043, 19.273626, 19.276686, 19.290142, 19.277807, 19.276081, 19.284689, 19.289917, 19.290003, 19.284868, 19.275778, 19.270035, 19.27149, 19.27132, 19.271524, 19.27438, 19.26817, 19.261402, 19.257446, 19.259716, 19.251305, 19.25465, 19.249798, 19.24574, 19.245998, 19.251587, 19.252472, 19.25991, 19.249537, 19.246084, 19.24335, 19.23914, 19.241203, 19.24003, 19.244768, 19.2486, 19.245455, 19.250608, 19.251448, 19.235973, 19.226868, 19.223612, 19.223743, 19.229542, 19.22866, 19.224974, 19.224123, 19.22584, 19.219652, 19.219387, 19.217928, 19.219084, 19.218153, 19.221548, 19.224339, 19.224092, 19.223335, 19.224087, 19.224789, 19.22732, 19.226864, 19.228405, 19.229921, 19.232183, 19.230883, 19.231564, 19.23449, 19.232323, 19.232635, 19.232767, 19.235292, 19.234924, 19.23751, 19.2368, 19.235548, 19.236855, 19.23604, 19.237398, 19.237244, 19.238392, 19.24372, 19.24148, 19.244251, 19.24296, 19.243093, 19.241936, 19.246796, 19.246525, 19.24805, 19.250214, 19.251919, 19.253353, 19.255644, 19.254763, 19.255602, 19.258553, 19.267473, 19.262396, 19.264572, 19.262718, 19.268805, 19.270445, 19.271393, 19.276188, 19.27527, 19.280876, 19.280005, 19.282377, 19.287985, 19.285114, 19.291264, 19.288721, 19.289547, 19.292873, 19.295918, 19.299725, 19.300909, 19.301996, 19.304144, 19.307343, 19.307337, 19.309685, 19.312494, 19.31371, 19.318758, 19.318768, 19.320065, 19.323029, 19.322807, 19.32767, 19.327637, 19.330345, 19.332201, 19.334112, 19.3356, 19.338406, 19.339657, 19.345337, 19.344332, 19.345486, 19.34843, 19.351723, 19.354471, 19.353369, 19.35179, 19.351501, 19.3496, 19.346682, 19.349928, 19.344347, 19.344938, 19.345446, 19.345804, 19.343779, 19.342302, 19.341963, 19.345158, 19.347076, 19.344942, 19.342737, 19.351748, 19.34961, 19.344292, 19.354958, 19.35861, 19.35946, 19.359348, 19.35864, 19.363293, 19.366442, 19.36853, 19.373234, 19.372192, 19.372679, 19.37294, 19.373941, 19.376152, 19.371761, 19.371454, 19.373695, 19.370993, 19.369274, 19.373064, 19.375296, 19.375547, 19.373474, 19.371838, 19.36932, 19.370586, 19.371243, 19.375235, 19.372177, 19.368504, 19.3747, 19.368073, 19.365904, 19.36918, 19.370079, 19.37505, 19.374321, 19.379097, 19.381538, 19.38279, 19.385387, 19.391785, 19.393473, 19.390923, 19.395279, 19.397089, 19.397818, 19.397223, 19.402744, 19.405813, 19.409164, 19.412525, 19.41328, 19.41619, 19.418736, 19.421516, 19.421522, 19.42052, 19.421907, 19.4187, 19.415539, 19.417965, 19.420004, 19.423647, 19.424257, 19.434647, 19.432922, 19.439781, 19.437742, 19.435541, 19.444956, 19.440613, 19.441248, 19.446856, 19.448175, 19.449602, 19.451748, 19.453966, 19.45646, 19.457602, 19.456373, 19.454823, 19.454449, 19.455208, 19.453781, 19.454094, 19.454243, 19.455574, 19.455748, 19.457565, 19.458588, 19.459742, 19.461334, 19.46346, 19.465288, 19.467018, 19.467825, 19.471174, 19.472298, 19.477238, 19.479343, 19.48127, 19.483238, 19.484959, 19.488354, 19.490984, 19.495708, 19.495205, 19.500137, 19.503256, 19.507011, 19.510643, 19.509975, 19.515093, 19.520374, 19.51741, 19.518745, 19.52056, 19.520334, 19.520844, 19.520575, 19.522959, 19.519852, 19.51777, 19.51591, 19.520061, 19.522955, 19.516983, 19.519312, 19.521059, 19.520884, 19.5193, 19.515776, 19.513968, 19.522287, 19.516357, 19.520956, 19.520777, 19.527369, 19.52337, 19.526022, 19.533262, 19.525597, 19.527205, 19.529743, 19.527311, 19.53334, 19.537468, 19.54071, 19.548538, 19.549232, 19.541286, 19.55047, 19.542822, 19.546005, 19.549623, 19.548868, 19.551514, 19.55175, 19.556793, 19.55669, 19.559698, 19.563976, 19.570284, 19.563616, 19.562254, 19.565702, 19.565481, 19.572777, 19.566912, 19.570906, 19.576212, 19.579226, 19.577658, 19.577374, 19.587082, 19.5864, 19.580177, 19.581549, 19.586723, 19.586851, 19.591387, 19.593506, 19.598639, 19.598654, 19.59551, 19.600027, 19.595486, 19.59883, 19.606575, 19.61232, 19.609516, 19.608606, 19.611074, 19.61941, 19.626905, 19.615648, 19.621832, 19.626688, 19.62135, 19.630856, 19.630362, 19.631073, 19.638033, 19.636892, 19.641136, 19.639624, 19.642443, 19.643385, 19.641933, 19.644312, 19.652819, 19.656101, 19.66162, 19.660852, 19.673164, 19.669056, 19.668577, 19.672567, 19.675507, 19.673658, 19.671486, 19.677431, 19.668995, 19.680603, 19.6814, 19.682987, 19.68209, 19.685335, 19.682755, 19.69005, 19.692059, 19.688414, 19.69075, 19.693495, 19.695076, 19.696667, 19.695797, 19.699097, 19.697603, 19.699148, 19.70571, 19.705713, 19.702177, 19.700684, 19.697182, 19.698727, 19.700312, 19.702244, 19.702969, 19.702995, 19.706924, 19.71038, 19.707846, 19.710978, 19.71145, 19.71487, 19.714098, 19.716066, 19.71653, 19.718084, 19.720798, 19.719208, 19.720964, 19.721355, 19.722546, 19.723173, 19.726624, 19.727362, 19.72731, 19.728567, 19.728289, 19.728664, 19.730467, 19.732805, 19.733574, 19.735052, 19.73431, 19.734728, 19.735758, 19.736206, 19.736382, 19.735937, 19.735746, 19.736406, 19.734692, 19.735437, 19.73397, 19.734325, 19.73411, 19.733908, 19.73445, 19.732857, 19.733316, 19.732862, 19.734346, 19.732254, 19.732084, 19.733223, 19.73275, 19.733053, 19.732353, 19.732388, 19.732975, 19.732584, 19.733644, 19.735788, 19.736391, 19.736675, 19.736525, 19.735022, 19.735092, 19.736282, 19.736467, 19.73689, 19.737658, 19.738317, 19.738586, 19.739147, 19.740198, 19.740343, 19.741192, 19.743557, 19.743397, 19.742975, 19.743093, 19.742697, 19.743757, 19.744062, 19.744598, 19.745304, 19.745329, 19.745686, 19.746216, 19.74657, 19.747478, 19.748848, 19.748745, 19.749481, 19.749905, 19.752213, 19.752254, 19.752197, 19.751064, 19.752146, 19.752249, 19.752909, 19.75257, 19.753403, 19.7533, 19.753466, 19.753708, 19.754608, 19.754635, 19.754063, 19.75445, 19.755331, 19.756655, 19.756407, 19.757402, 19.755783, 19.755074, 19.755268, 19.753506, 19.753378, 19.752691, 19.752533, 19.751755, 19.751137, 19.750616, 19.750513, 19.74974, 19.749502, 19.749868, 19.749704, 19.749462, 19.749271, 19.749744, 19.74956, 19.749605, 19.749895, 19.750565, 19.750898, 19.751007, 19.750677, 19.7518, 19.75164, 19.752104, 19.752522, 19.75195, 19.752228, 19.753496, 19.753021, 19.75412, 19.753521, 19.752842, 19.753218, 19.75348, 19.754593, 19.754208, 19.754417, 19.755331, 19.754711, 19.758036, 19.755077, 19.755625, 19.756433, 19.756334, 19.755753, 19.755465, 19.754381, 19.754692, 19.754738, 19.755402, 19.755217, 19.756128, 19.755589, 19.75548, 19.75564, 19.755552, 19.755589, 19.755228, 19.754568, 19.754501, 19.754423, 19.754196, 19.76461, 19.756525, 19.758566, 19.760168, 19.757679, 19.760406, 19.759148, 19.761518, 19.757463, 19.756021, 19.755737, 19.75548, 19.75601, 19.755573, 19.75548, 19.755383, 19.756613, 19.75704, 19.756021, 19.75647, 19.756077, 19.756319, 19.757164, 19.756386, 19.757294, 19.756603, 19.756212, 19.756573, 19.757767, 19.760529, 19.764065, 19.759138, 19.759571, 19.758417, 19.75799, 19.759607, 19.758932, 19.757542, 19.757118, 19.757727, 19.760046, 19.754614, 19.754347, 19.75684, 19.760319, 19.772026, 19.773615, 19.772995, 19.766321, 19.762066, 19.776604, 19.768532, 19.76458, 19.765194, 19.76279, 19.78236, 19.783386, 19.763926, 19.766075, 19.76375, 19.769985, 19.781557, 19.772676, 19.770742, 19.775005, 19.774805, 19.778221, 19.79734, 19.773727, 19.77865, 19.777386, 19.781918, 19.802893, 19.789066, 19.788979, 19.79268, 19.80083, 19.799965, 19.793634, 19.793484, 19.796495, 19.79946, 19.797186, 19.79962, 19.805244, 19.80297, 19.802382, 19.807224, 19.80477, 19.807858, 19.811535, 19.816113, 19.817614, 19.81946, 19.820692, 19.822475, 19.822502, 19.823383, 19.822853, 19.820925, 19.821428, 19.821712, 19.819185, 19.819784, 19.81804, 19.816195, 19.814112, 19.811152, 19.811033, 19.813591, 19.81301, 19.81011, 19.807688, 19.807116, 19.808487, 19.803898, 19.80301, 19.800419, 19.798237, 19.797386, 19.792175, 19.791325, 19.79021, 19.787031, 19.78404, 19.78338, 19.779943, 19.77902, 19.776897, 19.775, 19.775135, 19.775, 19.774733, 19.773912, 19.771887, 19.769176, 19.766745, 19.76558, 19.766363, 19.76627, 19.762636, 19.762436, 19.766106, 19.767656, 19.76809, 19.768496, 19.767786, 19.762445, 19.763435, 19.763926, 19.761915, 19.760468, 19.760477, 19.758596, 19.756649, 19.755253, 19.753517, 19.75714, 19.753305, 19.755068, 19.755701, 19.755453, 19.754686, 19.763863, 19.77163, 19.762596, 19.76425, 19.776798, 19.764853, 19.770945, 19.772991, 19.779135, 19.779531, 19.77633, 19.773897, 19.780603, 19.78064, 19.779078, 19.78684, 19.779392, 19.781185, 19.78167, 19.781366, 19.781385, 19.781715, 19.779762, 19.77865, 19.778221, 19.777536, 19.77602, 19.775866, 19.775175, 19.77366, 19.772825, 19.772856, 19.772789, 19.772526, 19.77231, 19.772774, 19.77565, 19.774563, 19.773794, 19.774635, 19.777128, 19.778572, 19.777454, 19.779108, 19.780952, 19.784382, 19.78403, 19.785252, 19.78917, 19.789005, 19.78781, 19.79088, 19.790396, 19.790655, 19.795336, 19.79134, 19.79082, 19.791464, 19.790026, 19.792793, 19.79038, 19.795948, 19.794561, 19.79214, 19.805738, 19.798216, 19.800413, 19.79497, 19.794846, 19.798721, 19.80532, 19.800068, 19.796432, 19.794954, 19.794743, 19.79197, 19.797083, 19.798124, 19.793371, 19.795351, 19.790783, 19.803331, 19.801443, 19.797985, 19.796516, 19.800434, 19.795391, 19.802729, 19.801186, 19.80777, 19.8109, 19.808771, 19.811117, 19.816278, 19.819794, 19.82097, 19.82621, 19.828499, 19.825184, 19.83443, 19.829836, 19.829933, 19.828773, 19.82968, 19.830753, 19.830273, 19.828949, 19.829903, 19.829845, 19.829155, 19.83605, 19.8341, 19.833496, 19.83158, 19.8303, 19.827246, 19.828695, 19.823147, 19.819118, 19.82114, 19.829506, 19.822977, 19.82475, 19.825384, 19.827112, 19.824528, 19.829428, 19.83161, 19.838114, 19.84114, 19.838108, 19.845901, 19.837458, 19.84505, 19.853664, 19.846552, 19.8468, 19.839367, 19.837706, 19.839996, 19.839237, 19.838516, 19.836246, 19.83948, 19.839867, 19.840242, 19.838387, 19.842894, 19.837706, 19.840351, 19.842157, 19.839125, 19.844303, 19.84476, 19.838526, 19.84424, 19.83917, 19.836353, 19.834982, 19.83805, 19.8341, 19.836988, 19.837376, 19.837633, 19.836143, 19.842615, 19.842642, 19.84374, 19.841068, 19.848465, 19.853401, 19.850048, 19.85106, 19.853134, 19.852148, 19.851818, 19.85123, 19.851494, 19.851658, 19.850002, 19.86807, 19.850178, 19.850922, 19.846752, 19.847826, 19.84828, 19.847466, 19.846437, 19.845303, 19.845684, 19.843735, 19.84571, 19.84293, 19.843765, 19.841465, 19.841383, 19.84341, 19.84467, 19.845335, 19.848946, 19.853222, 19.849941, 19.852804, 19.86109, 19.85948, 19.864473, 19.85922, 19.86581, 19.862017, 19.86891, 19.862455, 19.862198, 19.86096, 19.86049, 19.859665, 19.85965, 19.858938, 19.861795, 19.859407, 19.859783, 19.859919, 19.860739, 19.858845, 19.862167, 19.863829, 19.863714, 19.862724, 19.866388, 19.865768, 19.86842, 19.8634, 19.863705, 19.865236, 19.86582, 19.865656, 19.874323, 19.868921, 19.872347, 19.878286, 19.883318, 19.883757, 19.884438, 19.886316, 19.891142, 19.883411, 19.890062, 19.8968, 19.897713, 19.900251, 19.89829, 19.894781, 19.89829, 19.895765, 19.900045, 19.896328, 19.899576, 19.89875, 19.896969, 19.897955, 19.896835, 19.899622, 19.904577, 19.916967, 19.909166, 19.909124, 19.911236, 19.910963, 19.911459, 19.91437, 19.91599, 19.913347, 19.922253, 19.918293, 19.91532, 19.918505, 19.925104, 19.92656, 19.921593, 19.923214, 19.927675, 19.92897, 19.931015, 19.943083, 19.94017, 19.94095, 19.946527, 19.951683, 19.954466, 19.953201, 19.956388, 19.963537, 19.973156, 19.966383, 19.971798, 19.963713, 19.966295, 19.972406, 19.968536, 19.97638, 19.974556, 19.97686, 19.98103, 19.980755, 19.979527, 19.986998, 19.986042, 19.992144, 19.98692, 19.986166, 19.986336, 19.989798, 19.99309, 19.988703, 19.992878, 19.991177, 19.990946, 19.999704, 19.99345, 19.995493, 19.995424, 20.00218, 19.999187, 20.000355, 19.999777, 20.001001, 19.999989, 20.002014, 20.00602, 20.002686, 20.007595, 20.016657, 20.01572, 20.012867, 20.024374, 20.020182, 20.021267, 20.019598, 20.021914, 20.021412, 20.022823, 20.023703, 20.022854, 20.02123, 20.022596, 20.024529, 20.023252, 20.022978, 20.023428, 20.026121, 20.027548, 20.031006, 20.029352, 20.030561, 20.033058, 20.033628, 20.043322, 20.04418, 20.048203, 20.048311, 20.043509, 20.04097, 20.045975, 20.045452, 20.045137, 20.04418, 20.04568, 20.04508, 20.045788, 20.043213, 20.043802, 20.043766, 20.04067, 20.039103, 20.035091, 20.034714, 20.03387, 20.033792, 20.033209, 20.03095, 20.036264, 20.035292, 20.034817, 20.037355, 20.037685, 20.03857, 20.040897, 20.042841, 20.040834, 20.039455, 20.036053, 20.034487, 20.033943, 20.034067, 20.030428, 20.031942, 20.034155, 20.033587, 20.032284, 20.035826, 20.034222, 20.037706, 20.037878, 20.040907, 20.04051, 20.043911, 20.043255, 20.041533, 20.041653, 20.037086, 20.039547, 20.046125, 20.040995, 20.03815, 20.034233, 20.035576, 20.037186, 20.032604, 20.030785, 20.030537, 20.027802, 20.033173, 20.03447, 20.043959, 20.03978, 20.046642, 20.043518, 20.040958, 20.043533, 20.043684, 20.043493, 20.043524, 20.042913, 20.044004, 20.04448, 20.039598, 20.044355, 20.042889, 20.043425, 20.041248, 20.043224, 20.03962, 20.04055, 20.039656, 20.038317, 20.031002, 20.026731, 20.021385, 20.014647, 20.010098, 20.000603, 20.001328, 19.999239, 19.993834, 19.997126, 20.004562, 20.00663, 20.011694, 20.008749, 20.013344, 20.013363, 20.01891, 20.014997, 20.00771, 19.998423, 19.994066, 19.989204, 19.992403, 19.984709, 19.985065, 19.98788, 19.989447, 19.985725, 19.98323, 19.976797, 19.973068, 19.971172, 19.979427, 19.974586, 19.971336, 19.964048, 19.96005, 19.95973, 19.959373, 19.956512, 19.956491, 19.95256, 19.946436, 19.943027, 19.939014, 19.934278, 19.931227, 19.935204, 19.927086, 19.924128, 19.927996, 19.924593, 19.924835, 19.923565, 19.925192, 19.92309, 19.921738, 19.924034, 19.923492, 19.927654, 19.927996, 19.929348, 19.9323, 19.936737, 19.936008, 19.939644, 19.94568, 19.943115, 19.942692, 19.944075, 19.944933, 19.945045, 19.946182, 19.94925, 19.95116, 19.948868, 19.949875, 19.949854, 19.949802, 19.94859, 19.944918, 19.944876, 19.944386, 19.944147, 19.94265, 19.942123, 19.943161, 19.940294, 19.939798, 19.939169, 19.938818, 19.938648, 19.938261, 19.936855, 19.93146, 19.927158, 19.926725, 19.920591, 19.919455, 19.919104, 19.918411, 19.917746, 19.91644, 19.914364, 19.913342, 19.912537, 19.909895, 19.909542, 19.90854, 19.907757, 19.90594, 19.904339, 19.901144, 19.900194, 19.900076, 19.899426, 19.897964, 19.896524, 19.89446, 19.894373, 19.89623, 19.893867, 19.895317, 19.893835, 19.891296, 19.890516, 19.889227, 19.891394, 19.890131, 19.88885, 19.887463, 19.884396, 19.88485, 19.884928, 19.88385, 19.882023, 19.880924, 19.877306, 19.87616, 19.874292, 19.87082, 19.870722, 19.870691, 19.869886, 19.866806, 19.867311, 19.863974, 19.863947, 19.863312, 19.864313, 19.863241, 19.861961, 19.863611, 19.86132, 19.859795, 19.858288, 19.857008, 19.85735, 19.858545, 19.85512, 19.859026, 19.854832, 19.85413, 19.858082, 19.860073, 19.858143, 19.856373, 19.856688, 19.85673, 19.865934, 19.85413, 19.855274, 19.858839, 19.861507, 19.856838, 19.854975, 19.863039, 19.86011, 19.857147, 19.86066, 19.856808, 19.865923, 19.864706, 19.872765, 19.871202, 19.871588, 19.870607, 19.869778, 19.865953, 19.878017, 19.878674, 19.88645, 19.891127, 19.899858, 19.897774, 19.905548, 19.90067, 19.901299, 19.906786, 19.911547, 19.908289, 19.914309, 19.913889, 19.915583, 19.921091, 19.925419, 19.941813, 19.954487, 19.961218, 19.980099, 19.982956, 19.970345, 19.980146, 19.98766, 19.992065, 19.983473, 19.97669, 19.989136, 19.99295, 19.993824, 20.009626, 20.01049, 20.013468, 20.013172, 20.005766, 20.002577, 20.007307, 20.000944, 19.99821, 19.986387, 19.980522, 20.00788, 20.026592, 20.009073, 20.01322, 20.037579, 19.998459, 20.041565, 20.10723, 20.043436, 20.049765, 20.043095, 20.0789, 20.080347, 20.056002, 20.046564, 20.10158, 20.093819, 20.08109, 20.16835, 20.06833, 20.084568, 20.049221, 20.062853, 20.06649, 20.080673, 20.121239, 20.097227, 20.07503, 20.083658, 20.102257, 20.10263, 20.070927, 20.083967, 20.081738, 20.09981, 20.116732, 20.12244, 20.086668, 20.04868, 20.036833, 20.013002, 19.998444, 19.987839, 19.995085, 20.018993, 20.014465, 20.014475, 20.007673, 20.004923, 20.01784, 20.02672, 20.035397, 20.062471, 20.071217, 20.067348, 20.06003, 20.072552, 20.10126, 20.091915, 20.091, 20.100307, 20.096363, 20.146675, 20.120852, 20.097782, 20.077211, 20.06368, 20.051994, 20.053793, 20.056038, 20.08926, 20.117384, 20.0717, 20.042944, 20.047567, 20.040245, 20.022358, 19.978674, 19.982336, 20.000841, 19.990738, 19.987246, 19.996775, 19.968197, 19.947622, 19.950096, 19.922909, 19.931036, 19.915686, 19.91109, 19.907787, 19.912739, 19.882244, 19.91135, 19.889717, 19.895395, 19.886827, 19.862782, 19.849394, 19.846912, 19.840992, 19.843178, 19.831491, 19.82855, 19.840094, 19.834837, 19.832884, 19.818562, 19.812456, 19.812183, 19.818676, 19.82553, 19.82295, 19.82098, 19.806341, 19.794092, 19.796278, 19.794067, 19.784695, 19.782597, 19.784561, 19.77436, 19.763374, 19.757963, 19.755835, 19.763332, 19.756195, 19.749023, 19.742197, 19.740955, 19.739405, 19.73096, 19.724709, 19.72293, 19.71893, 19.719347, 19.71325, 19.715483, 19.715628, 19.727634, 19.742275, 19.730373, 19.727346, 19.729364, 19.738024, 19.729937, 19.72817, 19.726702, 19.72923, 19.73087, 19.736664, 19.731667, 19.734495, 19.733208, 19.739931, 19.749817, 19.755783, 19.753717, 19.765461, 19.764492, 19.765915, 19.778078, 19.771908, 19.777346, 19.7737, 19.772207, 19.773443, 19.777748, 19.77645, 19.78402, 19.776104, 19.773022, 19.76623, 19.777288, 19.758963, 19.779432, 19.79005, 19.798212, 19.796532, 19.789618, 19.780005, 19.77228, 19.76259, 19.757933, 19.756052, 19.756067, 19.768068, 19.772392, 19.770552, 19.768295, 19.744799, 19.743654, 19.752981, 19.760246, 19.76391, 19.773006, 19.760298, 19.740828, 19.733553, 19.725145, 19.719692, 19.708197, 19.7294, 19.722843, 19.725702, 19.714767, 19.71676, 19.70983, 19.725254, 19.704838, 19.705235, 19.71485, 19.725863, 19.74094, 19.744377, 19.763441, 19.763632, 19.760683, 19.776707, 19.770018, 19.784298, 19.783123, 19.76947, 19.770517, 19.761467, 19.764435, 19.773212, 19.77294, 19.776165, 19.780449, 19.77569, 19.77616, 19.769176, 19.774305, 19.760906, 19.754887, 19.755196, 19.773186, 19.754166, 19.750471, 19.746376, 19.752172, 19.738977, 19.745644, 19.731842, 19.726469, 19.714643, 19.717539, 19.712759, 19.710056, 19.707203, 19.705095, 19.698536, 19.690468, 19.684547, 19.688053, 19.680082, 19.683512, 19.684088, 19.678503, 19.679249, 19.673, 19.685545, 19.680948, 19.679893, 19.678064, 19.665634, 19.664341, 19.65499, 19.655983, 19.654377, 19.658417, 19.654476, 19.651546, 19.670513, 19.670504, 19.664831, 19.667095, 19.657965, 19.656452, 19.663147, 19.659813, 19.656189, 19.656622, 19.657337, 19.655807, 19.66689, 19.666092, 19.658998, 19.669804, 19.656647, 19.665464, 19.659971, 19.670174, 19.662071, 19.673325, 19.672907, 19.66671, 19.663713, 19.65762, 19.679876, 19.667667, 19.680304, 19.676943, 19.68881, 19.676325, 19.677443, 19.681776, 19.692522, 19.68761, 19.67911, 19.675137, 19.681112, 19.68501, 19.690601, 19.682121, 19.694613, 19.698896, 19.693104, 19.70487, 19.69576, 19.689531, 19.702408, 19.691807, 19.688414, 19.681479, 19.680124, 19.689062, 19.689062, 19.687254, 19.689808, 19.697815, 19.701008, 19.734196, 19.714588, 19.726408, 19.72018, 19.726902, 19.73614, 19.74448, 19.727726, 19.72771, 19.735628, 19.744205, 19.740137, 19.73225, 19.738863, 19.742727, 19.752615, 19.747467, 19.746216, 19.75262, 19.751234, 19.778706, 19.76829, 19.779556, 19.766775, 19.771248, 19.774563, 19.792814, 19.792685, 19.800186, 19.796305, 19.805475, 19.84229, 19.812147, 19.811142, 19.80332, 19.790495, 19.78452, 19.790861, 19.817005, 19.790014, 19.818819, 19.816902, 19.825287, 19.828505, 19.833517, 19.835411, 19.849709, 19.839815, 19.842224, 19.857983, 19.861631, 19.842306, 19.843513, 19.862349, 19.85623, 19.852205, 19.855852, 19.85022, 19.884045, 19.866652, 19.852262, 19.879452, 19.87693, 19.892107, 19.89034, 19.900696, 19.891384, 19.891079, 19.90355, 19.906694, 19.934904, 19.917793, 19.919027, 19.91217, 19.9323, 19.937466, 19.936768, 19.92583, 19.954859, 19.944994, 19.951487, 19.946053, 19.956713, 19.933613, 19.934732, 19.931662, 19.929264, 19.939386, 19.944649, 19.938374, 19.922192, 19.931583, 19.930622, 19.961874, 19.93041, 19.92518, 19.934006, 19.970707, 19.9434, 19.934254, 19.926968, 19.921118, 19.912067, 19.839764, 19.801563, 19.819675, 19.806528, 19.742636, 19.7462, 19.746834, 19.69696, 19.722643, 19.69002, 19.636017, 19.628674, 19.618488, 19.589464, 19.532179, 19.527641, 19.49636, 19.487238, 19.482452, 19.47089, 19.45951, 19.451902, 19.44204, 19.437614, 19.427856, 19.435818, 19.43472, 19.44319, 19.446491, 19.454828, 19.456585, 19.45223, 19.464144, 19.459122, 19.455265, 19.464384, 19.474861, 19.4718, 19.474224, 19.472437, 19.488373, 19.487228, 19.494959, 19.49123, 19.52723, 19.53074, 19.506456, 19.505522, 19.51424, 19.507685, 19.525715, 19.542181, 19.527193, 19.536613, 19.542961, 19.559795, 19.561005, 19.556902, 19.570515, 19.592411, 19.607985, 19.597044, 19.607494, 19.63452, 19.649937, 19.657825, 19.684423, 19.689138, 19.69856, 19.704185, 19.72406, 19.728128, 19.715294, 19.739704, 19.767769, 19.785887, 19.824333, 19.805124, 19.819908, 19.852148, 19.842194, 19.858067, 19.853437, 19.874752, 19.878637, 19.881687, 19.903343, 19.871475, 19.893583, 19.91088, 19.892633, 19.888622, 19.893051, 19.90949, 19.902729, 19.891178, 19.90994, 19.888391, 19.894258, 19.902575, 19.89925, 19.915552, 19.890718, 19.870398, 19.880356, 19.92544, 19.884861, 19.878323, 19.876965, 19.877466, 19.86827, 19.843235, 19.833399, 19.857952, 19.831387, 19.829494, 19.817572, 19.836504, 19.811275, 19.811596, 19.818573, 19.787598, 19.813555, 19.869923, 19.789526, 19.749838, 19.705456, 19.69001, 19.694649, 19.685448, 19.685406, 19.711487, 19.70053, 19.682055, 19.66185, 19.656853, 19.682976, 19.63437, 19.62516, 19.610731, 19.60498, 19.561348, 19.54878, 19.558628, 19.620525, 19.5922, 19.585915, 19.583813, 19.599209, 19.601858, 19.626503, 19.63349, 19.621456, 19.59856, 19.591808, 19.582985, 19.573368, 19.614141, 19.592405, 19.613796, 19.60569, 19.612562, 19.628607, 19.622465, 19.621601, 19.591274, 19.564772, 19.564695, 19.571291, 19.563148, 19.574938, 19.584517, 19.576397, 19.611856, 19.598433, 19.634035, 19.64091, 19.657553, 19.658089, 19.638512, 19.640081, 19.666473, 19.654459, 19.686008, 19.65795, 19.69311, 19.674385, 19.720072, 19.694052, 19.716833, 19.734196, 19.725914, 19.755438, 19.75564, 19.775671, 19.756495, 19.768377, 19.749002, 19.753923, 19.76827, 19.78819, 19.787891, 19.771908, 19.80035, 19.77901, 19.792727, 19.81409, 19.791386, 19.813591, 19.819294, 19.816587, 19.814907, 19.830284, 19.833496, 19.873251, 19.842781, 19.881966, 19.919119, 19.945469, 19.951088, 20.001125, 19.973032, 19.979769, 19.966358, 20.078356, 20.04962, 20.070524, 20.072153, 20.145868, 20.185757, 20.240732, 20.180075, 20.200521, 20.233166, 20.203043, 20.21695, 20.257755, 20.325455, 20.31758, 20.316967, 20.307266, 20.322279, 20.385672, 20.342335, 20.388798, 20.384695, 20.374706, 20.379322, 20.415659, 20.431759, 20.433031, 20.412994, 20.408527, 20.394402, 20.407837, 20.369238, 20.353935, 20.338724, 20.339424, 20.332745, 20.32049, 20.270117, 20.217836, 20.184359, 20.154686, 20.008314, 19.96836, 19.934961, 19.877512, 19.838789, 19.797907, 19.768183, 19.68745, 19.694555, 19.644215, 19.647058, 19.594355, 19.551992, 19.559292, 19.526741, 19.507088, 19.494152, 19.476273, 19.456476, 19.44555, 19.401466, 19.383509, 19.376984, 19.363949, 19.353184, 19.352615, 19.35499, 19.35961, 19.36694, 19.355415, 19.364437, 19.373674, 19.403458, 19.385458, 19.38218, 19.38142, 19.367987, 19.354082, 19.345722, 19.33785, 19.354462, 19.369387, 19.388777, 19.488256, 19.422697, 19.453405, 19.451836, 19.465807, 19.462479, 19.46328, 19.485199, 19.480793, 19.479118, 19.478542, 19.489227, 19.463522, 19.47595, 19.449581, 19.463692, 19.485168, 19.467367, 19.446604, 19.464745, 19.445639, 19.442762, 19.461704, 19.44242, 19.468605, 19.552692, 19.500692, 19.487978, 19.522861, 19.495165, 19.54193, 19.508522, 19.537344, 19.562145, 19.507263, 19.593485, 19.552938, 19.548801, 19.563698, 19.573893, 19.531075, 19.58065, 19.603695, 19.56743, 19.632301, 19.581375, 19.7049, 19.58391, 19.655962, 19.64197, 19.656374, 19.70042, 19.610407, 19.677958, 19.673452, 19.650625, 19.612686, 19.851406, 19.637072, 19.694113, 19.707409, 19.729952, 19.718542, 19.67254, 19.684464, 19.722834, 19.723745, 19.667322, 19.781542, 19.684748, 19.811415, 19.744804, 19.732327, 19.69799, 19.70109, 19.68572, 19.662237, 19.740328, 19.672104, 19.662756, 19.690432, 19.642315, 19.627893, 19.624826, 19.627321, 19.634647, 19.612556, 19.640005, 19.613087, 19.610561, 19.606857, 19.613132, 19.59674, 19.611004, 19.590805, 19.573538, 19.589952, 19.582361, 19.585915, 19.591942, 19.615324, 19.600325, 19.603956, 19.571148, 19.56213, 19.586845, 19.549093, 19.576536, 19.598408, 19.57362, 19.541945, 19.546122, 19.548765, 19.551868, 19.54695, 19.552002, 19.557575, 19.541908, 19.54088, 19.531696, 19.534399, 19.530832, 19.52422, 19.520504, 19.527302, 19.536259, 19.52721, 19.520267, 19.51855, 19.51422, 19.512653, 19.51054, 19.505444, 19.498129, 19.496798, 19.49421, 19.492268, 19.494862, 19.49089, 19.48603, 19.479729, 19.477407, 19.463512, 19.457981, 19.440355, 19.428959, 19.441244, 19.437538, 19.406609, 19.402985, 19.399086, 19.397732, 19.40047, 19.401442, 19.397161, 19.397408, 19.389301, 19.39218, 19.394007, 19.39398, 19.39157, 19.391256, 19.394909, 19.406715, 19.402908, 19.41467, 19.416939, 19.415764, 19.416441, 19.41757, 19.423006, 19.437254, 19.44168, 19.444504, 19.439663, 19.434565, 19.441618, 19.455177, 19.447866, 19.44996, 19.46134, 19.455608, 19.462627, 19.461786, 19.468632, 19.47859, 19.494728, 19.484692, 19.475985, 19.491394, 19.493433, 19.498318, 19.504103, 19.486397, 19.503004, 19.50756, 19.521942, 19.507385, 19.510818, 19.522066, 19.522497, 19.518654, 19.513695, 19.523037, 19.537529, 19.542463, 19.52888, 19.534168, 19.575039, 19.571712, 19.575005, 19.57869, 19.596216, 19.576736, 19.571173, 19.584743, 19.586666, 19.578362, 19.59551, 19.5879, 19.608328, 19.617685, 19.60607, 19.607485, 19.604275, 19.61252, 19.629868, 19.631294, 19.645557, 19.6402, 19.664768, 19.698145, 19.697433, 19.713764, 19.720577, 19.719465, 19.70714, 19.714474, 19.756891, 19.735464, 19.734253, 19.758045, 19.776583, 19.773785, 19.786674, 19.818134, 19.819681, 19.789175, 19.852133, 19.80627, 19.864885, 19.885357, 19.893536, 19.958, 19.928719, 19.956516, 20.013287, 19.913677, 19.89991, 19.879917, 19.892237, 20.027626, 20.031265, 20.051481, 20.002966, 20.076803, 20.056772, 20.023117, 20.04813, 20.127476, 20.077036, 20.077139, 20.109446, 20.114826, 20.115469, 20.170956, 20.170412, 20.152437, 20.144594, 20.167227, 20.156404, 20.157558, 20.194864, 20.176409, 20.158419, 20.16936, 20.16793, 20.167812, 20.192999, 20.176134, 20.19505, 20.18959, 20.191797, 20.205261, 20.237259, 20.209318, 20.216578, 20.229029, 20.243677, 20.259813, 20.270802, 20.276474, 20.28812, 20.302235, 20.303204, 20.32695, 20.336285, 20.34491, 20.339907, 21.316433, 22.433838, 26.638023, 24.403727, 25.100468, 26.601774, 27.391539, 27.575779, 28.709026, 29.309935, 29.51387, 29.596525, 29.596876, 29.842253, 29.836094, 29.855976, 30.118168, 32.39682, 35.02877, 35.609524, 36.697197, 34.059414, 35.10359, 34.234417, 32.881092, 32.998287, 35.96515, 33.414772, 32.320404, 31.228168, 29.062532, 28.01052, 26.696669, 25.938372, 25.353086, 25.375103}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_REL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
DEPTH =
  {39.402702, 39.407234, 39.411766, 39.416298, 39.42083, 39.42536, 39.429893, 39.428757, 39.42762, 39.426483, 39.42535, 39.424213, 39.423077, 39.429874, 39.436676, 39.443474, 39.45027, 39.457073, 39.46387, 39.462734, 39.461594, 39.460457, 39.45932, 39.45818, 39.457043, 39.46669, 39.476334, 39.485977, 39.495625, 39.50527, 39.514915, 39.51773, 39.520546, 39.52336, 39.52618, 39.528996, 39.53181, 39.53749, 39.54317, 39.54885, 39.554527, 39.560207, 39.565887, 39.562485, 39.559086, 39.555683, 39.55228, 39.54888, 39.54548, 39.55001, 39.554543, 39.559074, 39.563602, 39.568134, 39.572666, 39.573235, 39.573807, 39.57438, 39.574947, 39.575516, 39.576088, 39.58458, 39.593067, 39.60156, 39.61005, 39.618538, 39.62703, 39.62364, 39.62025, 39.61686, 39.61347, 39.61008, 39.60669, 39.612347, 39.618004, 39.623665, 39.629322, 39.63498, 39.640636, 39.642906, 39.645176, 39.647446, 39.64971, 39.65198, 39.65425, 39.65708, 39.659912, 39.662743, 39.665577, 39.668407, 39.671238, 39.670113, 39.668983, 39.66786, 39.666733, 39.665604, 39.66448, 39.667885, 39.671288, 39.67469, 39.678097, 39.6815, 39.684906, 39.692265, 39.699627, 39.706985, 39.714344, 39.721706, 39.729065, 39.7302, 39.73134, 39.732475, 39.733612, 39.73475, 39.735886, 39.73135, 39.72681, 39.722275, 39.71774, 39.7132, 39.708664, 39.71263, 39.716595, 39.72056, 39.724525, 39.72849, 39.732456, 39.728493, 39.724525, 39.72056, 39.716595, 39.71263, 39.708664, 39.706394, 39.704124, 39.70185, 39.69958, 39.69731, 39.69504, 39.700153, 39.70526, 39.710373, 39.71548, 39.72059, 39.7257, 39.719475, 39.713245, 39.70702, 39.700794, 39.694565, 39.68834, 39.69343, 39.69852, 39.703613, 39.708706, 39.713795, 39.718887, 39.70585, 39.692806, 39.679768, 39.66673, 39.653687, 39.640648, 39.638947, 39.63725, 39.635548, 39.633846, 39.63215, 39.630447, 39.625916, 39.621387, 39.61686, 39.612328, 39.6078, 39.603268, 39.60157, 39.59987, 39.59817, 39.596474, 39.594772, 39.593075, 39.584003, 39.574936, 39.565865, 39.556793, 39.547726, 39.538654, 39.54206, 39.545467, 39.548874, 39.552277, 39.555683, 39.55909, 39.544933, 39.530777, 39.516617, 39.50246, 39.488304, 39.474148, 39.478664, 39.48318, 39.487698, 39.492214, 39.49673, 39.501247, 39.49445, 39.48765, 39.48085, 39.474052, 39.467255, 39.460457, 39.455925, 39.451393, 39.44686, 39.442326, 39.437794, 39.43326, 39.42873, 39.424202, 39.41967, 39.41514, 39.41061, 39.40608, 39.407787, 39.409492, 39.4112, 39.41291, 39.414616, 39.416325, 39.407818, 39.399307, 39.3908, 39.382294, 39.373783, 39.365276, 39.371513, 39.37775, 39.383987, 39.39023, 39.396465, 39.402702, 39.39703, 39.391357, 39.385685, 39.380013, 39.37434, 39.368668, 39.36812, 39.36757, 39.36702, 39.366474, 39.365925, 39.365376, 39.36763, 39.369884, 39.37214, 39.374397, 39.37665, 39.378906, 39.381737, 39.384567, 39.387398, 39.39023, 39.39306, 39.39589, 39.387966, 39.38004, 39.372116, 39.364193, 39.356266, 39.348343, 39.35173, 39.355118, 39.358505, 39.361893, 39.36528, 39.368668, 39.377182, 39.385696, 39.39421, 39.402725, 39.41124, 39.419754, 39.408985, 39.398212, 39.387444, 39.376675, 39.365902, 39.355133, 39.356262, 39.35739, 39.35852, 39.359646, 39.360775, 39.361904, 39.36926, 39.376614, 39.383972, 39.391327, 39.39868, 39.406036, 39.398113, 39.390186, 39.382263, 39.37434, 39.366413, 39.35849, 39.36642, 39.374355, 39.382286, 39.39022, 39.39815, 39.406086, 39.41516, 39.424236, 39.43331, 39.44239, 39.451466, 39.46054, 39.469032, 39.477524, 39.486015, 39.494503, 39.502995, 39.511486, 39.509792, 39.5081, 39.506405, 39.50471, 39.503017, 39.501324, 39.501312, 39.501297, 39.501286, 39.501274, 39.50126, 39.501247, 39.501255, 39.501263, 39.501274, 39.50128, 39.50129, 39.501297, 39.506954, 39.51261, 39.51827, 39.523926, 39.529583, 39.53524, 39.539223, 39.543205, 39.547188, 39.551167, 39.55515, 39.55913, 39.56479, 39.570446, 39.576103, 39.58176, 39.587418, 39.593075, 39.5976, 39.60212, 39.606644, 39.611168, 39.61569, 39.620213, 39.61966, 39.619106, 39.618553, 39.617996, 39.617443, 39.61689, 39.61518, 39.613472, 39.611763, 39.610054, 39.608345, 39.606636, 39.611744, 39.616856, 39.621964, 39.62707, 39.632183, 39.63729, 39.640682, 39.64407, 39.64746, 39.650852, 39.65424, 39.65763, 39.670673, 39.683716, 39.69676, 39.7098, 39.722843, 39.735886, 39.734173, 39.73246, 39.730743, 39.72903, 39.727318, 39.725605, 39.727318, 39.72903, 39.730743, 39.73246, 39.734173, 39.735886, 39.729633, 39.723385, 39.717133, 39.71088, 39.70463, 39.69838, 39.701786, 39.705193, 39.7086, 39.712006, 39.715412, 39.71882, 39.719967, 39.72111, 39.72226, 39.723408, 39.724552, 39.7257, 39.725693, 39.72569, 39.72568, 39.725674, 39.72567, 39.725662, 39.717728, 39.70979, 39.701855, 39.69392, 39.68598, 39.678047, 39.67975, 39.681446, 39.683147, 39.68485, 39.686546, 39.688248, 39.684845, 39.68144, 39.678036, 39.674633, 39.671227, 39.667824, 39.663307, 39.65879, 39.654274, 39.649754, 39.645237, 39.64072, 39.625984, 39.61125, 39.596516, 39.58178, 39.567047, 39.55231, 39.550613, 39.548916, 39.54722, 39.54552, 39.543823, 39.542126, 39.532475, 39.522823, 39.51317, 39.503517, 39.493866, 39.484215, 39.487625, 39.491035, 39.494446, 39.497856, 39.501266, 39.504677, 39.487118, 39.469555, 39.451996, 39.434437, 39.416874, 39.399315, 39.400444, 39.401573, 39.402702, 39.403828, 39.404957, 39.406086, 39.395885, 39.38568, 39.37548, 39.36528, 39.355076, 39.344875, 39.34658, 39.34828, 39.349987, 39.351692, 39.353394, 39.3551, 39.351692, 39.34829, 39.344883, 39.341476, 39.338074, 39.334667, 39.332417, 39.330166, 39.327915, 39.325665, 39.323414, 39.321163, 39.31605, 39.31094, 39.305824, 39.300713, 39.2956, 39.29049, 39.28596, 39.28143, 39.2769, 39.27237, 39.26784, 39.26331, 39.262737, 39.26217, 39.261597, 39.261024, 39.260456, 39.259884, 39.25819, 39.2565, 39.254807, 39.253117, 39.251427, 39.249733, 39.25312, 39.25651, 39.259903, 39.26329, 39.266678, 39.27007, 39.268936, 39.2678, 39.266666, 39.265533, 39.264397, 39.263264, 39.26838, 39.2735, 39.278614, 39.28373, 39.28885, 39.293964, 39.291687, 39.289413, 39.287136, 39.28486, 39.282585, 39.280308, 39.284855, 39.2894, 39.293945, 39.29849, 39.303032, 39.30758, 39.307564, 39.30755, 39.307533, 39.307518, 39.307503, 39.307487, 39.307495, 39.307503, 39.30751, 39.307518, 39.307526, 39.307533, 39.309788, 39.312042, 39.314297, 39.31655, 39.318806, 39.32106, 39.32957, 39.33808, 39.34659, 39.3551, 39.36361, 39.37212, 39.378353, 39.384586, 39.390816, 39.39705, 39.403282, 39.409515, 39.41064, 39.41177, 39.412895, 39.41402, 39.41515, 39.416275, 39.417416, 39.418552, 39.419693, 39.42083, 39.421967, 39.423107, 39.4265, 39.42989, 39.43328, 39.436676, 39.440067, 39.44346, 39.44686, 39.450264, 39.453667, 39.457073, 39.460476, 39.46388, 39.46332, 39.462765, 39.46221, 39.461655, 39.461098, 39.46054, 39.461098, 39.461655, 39.46221, 39.462765, 39.46332, 39.46388, 39.46897, 39.474064, 39.479156, 39.484253, 39.489346, 39.49444, 39.500114, 39.505787, 39.51146, 39.517136, 39.522808, 39.528484, 39.53074, 39.532993, 39.535248, 39.537502, 39.539757, 39.54201, 39.540325, 39.538643, 39.536957, 39.53527, 39.53359, 39.531902, 39.535854, 39.53981, 39.543762, 39.547714, 39.55167, 39.555622, 39.56469, 39.573757, 39.582825, 39.591892, 39.60096, 39.610027, 39.620228, 39.630432, 39.640633, 39.650833, 39.661037, 39.671238, 39.67408, 39.676918, 39.679756, 39.6826, 39.685436, 39.68828, 39.686012, 39.683743, 39.681473, 39.679207, 39.67694, 39.67467, 39.680336, 39.686, 39.691666, 39.697327, 39.70299, 39.708656, 39.711483, 39.714306, 39.717133, 39.719955, 39.72278, 39.725605, 39.72787, 39.73014, 39.732407, 39.734676, 39.736942, 39.739212, 39.732407, 39.7256, 39.718796, 39.71199, 39.705185, 39.69838, 39.70746, 39.716537, 39.725616, 39.73469, 39.74377, 39.75285, 39.746048, 39.739246, 39.732445, 39.725647, 39.718845, 39.712044, 39.709206, 39.706364, 39.703526, 39.700687, 39.697845, 39.695007, 39.688786, 39.682568, 39.676346, 39.670124, 39.663906, 39.657684, 39.653152, 39.648624, 39.644093, 39.63956, 39.635033, 39.6305, 39.6186, 39.606697, 39.594795, 39.582893, 39.57099, 39.55909, 39.56136, 39.563625, 39.565895, 39.56816, 39.570427, 39.572697, 39.56363, 39.55456, 39.545494, 39.53643, 39.527363, 39.518295, 39.513187, 39.508076, 39.502968, 39.49786, 39.49275, 39.48764, 39.474056, 39.460472, 39.44689, 39.433308, 39.419724, 39.40614, 39.395943, 39.385746, 39.37555, 39.365353, 39.355156, 39.34496, 39.340427, 39.335896, 39.331367, 39.326836, 39.322304, 39.317772, 39.313225, 39.308678, 39.30413, 39.299583, 39.295036, 39.29049, 39.28993, 39.289364, 39.288803, 39.288242, 39.287678, 39.287117, 39.277493, 39.267864, 39.25824, 39.248615, 39.238987, 39.229362, 39.22369, 39.218014, 39.21234, 39.20667, 39.200993, 39.19532, 39.19928, 39.20324, 39.2072, 39.211163, 39.215122, 39.21908, 39.215687, 39.21229, 39.208897, 39.2055, 39.202106, 39.19871, 39.19701, 39.19531, 39.193604, 39.191902, 39.1902, 39.1885, 39.186794, 39.18509, 39.183388, 39.181683, 39.179977, 39.178272, 39.17544, 39.17261, 39.16978, 39.16695, 39.16412, 39.16129, 39.17092, 39.180553, 39.190186, 39.199814, 39.209446, 39.219078, 39.217396, 39.215714, 39.214027, 39.212345, 39.210663, 39.20898, 39.215775, 39.222565, 39.229355, 39.23615, 39.24294, 39.249733, 39.249725, 39.24972, 39.249718, 39.24971, 39.249706, 39.2497, 39.255936, 39.262173, 39.26841, 39.274643, 39.28088, 39.287117, 39.285988, 39.284863, 39.283737, 39.282608, 39.281483, 39.280354, 39.28318, 39.286003, 39.288826, 39.291653, 39.294476, 39.297302, 39.306934, 39.316566, 39.326202, 39.335835, 39.345467, 39.3551, 39.36303, 39.370956, 39.378883, 39.386814, 39.39474, 39.40267, 39.403255, 39.40384, 39.404423, 39.405006, 39.40559, 39.406174, 39.41183, 39.41749, 39.423145, 39.428802, 39.43446, 39.440117, 39.437283, 39.43445, 39.43161, 39.428776, 39.42594, 39.423107, 39.42708, 39.43105, 39.43502, 39.438988, 39.44296, 39.44693, 39.445225, 39.443516, 39.44181, 39.440105, 39.438396, 39.43669, 39.446888, 39.457085, 39.467278, 39.477474, 39.48767, 39.497868, 39.49901, 39.50015, 39.50129, 39.502434, 39.503574, 39.504715, 39.502457, 39.500195, 39.497932, 39.495674, 39.493416, 39.491154, 39.49455, 39.49794, 39.501335, 39.50473, 39.50812, 39.511517, 39.51718, 39.522846, 39.52851, 39.53418, 39.539845, 39.54551, 39.556263, 39.567017, 39.577766, 39.58852, 39.599274, 39.610027, 39.61966, 39.62929, 39.638924, 39.64856, 39.65819, 39.667824, 39.671227, 39.674633, 39.678036, 39.68144, 39.684845, 39.688248, 39.688816, 39.689384, 39.689957, 39.690525, 39.691093, 39.69166, 39.69563, 39.699596, 39.70356, 39.707527, 39.711494, 39.71546, 39.72056, 39.72565, 39.730743, 39.73584, 39.740932, 39.74603, 39.756233, 39.766438, 39.77664, 39.78685, 39.797054, 39.80726, 39.80782, 39.808376, 39.808937, 39.809498, 39.810055, 39.810616, 39.811745, 39.812874, 39.814003, 39.815132, 39.81626, 39.81739, 39.812866, 39.808346, 39.80382, 39.799297, 39.794777, 39.790253, 39.78911, 39.787968, 39.786827, 39.785683, 39.784542, 39.783398, 39.77433, 39.765263, 39.756195, 39.747124, 39.738056, 39.72899, 39.72561, 39.722225, 39.718845, 39.715466, 39.712082, 39.708702, 39.70529, 39.701885, 39.698475, 39.695065, 39.691658, 39.688248, 39.67975, 39.671253, 39.662754, 39.654255, 39.64576, 39.63726, 39.625923, 39.614582, 39.60324, 39.591904, 39.580566, 39.569225, 39.566395, 39.56356, 39.56073, 39.5579, 39.555065, 39.552235, 39.537506, 39.52278, 39.508053, 39.493324, 39.4786, 39.46387, 39.45652, 39.449165, 39.44181, 39.43446, 39.42711, 39.419754, 39.412945, 39.406136, 39.399326, 39.392517, 39.385708, 39.3789, 39.373234, 39.36757, 39.3619, 39.356236, 39.35057, 39.344906, 39.334133, 39.32336, 39.312588, 39.301815, 39.291042, 39.28027, 39.275745, 39.271217, 39.266693, 39.26217, 39.25764, 39.253117, 39.251987, 39.250862, 39.249733, 39.248608, 39.247482, 39.246353, 39.24012, 39.233883, 39.227646, 39.221413, 39.21518, 39.208942, 39.202705, 39.196472, 39.190235, 39.184, 39.177765, 39.171528, 39.169827, 39.16813, 39.166428, 39.164726, 39.16303, 39.161327, 39.15849, 39.155647, 39.15281, 39.149967, 39.14713, 39.144287, 39.14996, 39.155632, 39.16131, 39.16698, 39.172653, 39.178326, 39.18399, 39.18966, 39.195324, 39.20099, 39.206657, 39.212322, 39.22082, 39.229317, 39.237816, 39.246315, 39.25481, 39.26331, 39.26106, 39.25881, 39.256554, 39.254303, 39.252052, 39.2498, 39.254887, 39.259968, 39.265053, 39.270138, 39.27522, 39.280304, 39.2837, 39.287094, 39.29049, 39.293888, 39.297283, 39.30068, 39.309185, 39.31769, 39.3262, 39.334705, 39.343212, 39.35172, 39.35569, 39.359657, 39.363625, 39.367596, 39.371563, 39.375534, 39.375538, 39.375546, 39.37555, 39.375557, 39.37556, 39.37557, 39.384632, 39.393692, 39.402756, 39.411816, 39.420876, 39.42994, 39.42483, 39.41972, 39.41461, 39.409504, 39.404392, 39.399284, 39.410065, 39.420845, 39.431625, 39.44241, 39.45319, 39.46397, 39.467915, 39.47186, 39.475807, 39.47975, 39.483696, 39.48764, 39.48595, 39.48426, 39.48257, 39.48088, 39.47919, 39.4775, 39.48203, 39.48656, 39.49109, 39.495617, 39.50015, 39.504677, 39.502975, 39.501274, 39.499573, 39.49787, 39.49617, 39.49447, 39.49447, 39.49447, 39.49447, 39.49447, 39.49447, 39.49447, 39.504105, 39.51374, 39.523376, 39.53301, 39.542645, 39.55228, 39.545483, 39.53868, 39.531883, 39.525085, 39.518284, 39.511486, 39.51488, 39.51828, 39.521675, 39.52507, 39.52847, 39.531864, 39.54659, 39.561314, 39.57604, 39.590763, 39.605488, 39.620213, 39.63157, 39.64292, 39.654274, 39.66563, 39.676983, 39.68834, 39.68834, 39.68834, 39.68834, 39.68834, 39.68834, 39.68834, 39.700222, 39.712105, 39.723988, 39.73587, 39.747753, 39.759636, 39.760757, 39.76188, 39.763, 39.76412, 39.76524, 39.76636, 39.77657, 39.786777, 39.79699, 39.807198, 39.817406, 39.827614, 39.82989, 39.83217, 39.834446, 39.836723, 39.839, 39.841278, 39.84977, 39.858257, 39.86675, 39.87524, 39.883728, 39.89222, 39.89505, 39.89788, 39.90071, 39.903545, 39.906376, 39.909206, 39.91544, 39.921677, 39.92791, 39.934143, 39.94038, 39.946613, 39.939816, 39.933014, 39.926216, 39.91942, 39.912617, 39.90582, 39.910343, 39.914867, 39.919395, 39.92392, 39.928444, 39.93297, 39.91994, 39.906914, 39.893883, 39.880856, 39.86783, 39.8548, 39.85196, 39.84912, 39.84628, 39.843437, 39.8406, 39.837757, 39.833805, 39.82985, 39.825897, 39.821945, 39.81799, 39.814037, 39.798172, 39.782307, 39.76644, 39.75058, 39.734715, 39.71885, 39.711487, 39.704124, 39.696762, 39.689396, 39.682034, 39.67467, 39.669003, 39.663338, 39.65767, 39.652, 39.646336, 39.640667, 39.628773, 39.616882, 39.60499, 39.593094, 39.581203, 39.56931, 39.56024, 39.551174, 39.542107, 39.533043, 39.523975, 39.514908, 39.504704, 39.4945, 39.4843, 39.474094, 39.46389, 39.453686, 39.445744, 39.4378, 39.429863, 39.42192, 39.41398, 39.406036, 39.399242, 39.39245, 39.38566, 39.378864, 39.37207, 39.365276, 39.35678, 39.348286, 39.33979, 39.331295, 39.3228, 39.314304, 39.305805, 39.297306, 39.288807, 39.280308, 39.27181, 39.26331, 39.264446, 39.265583, 39.266724, 39.26786, 39.268997, 39.270134, 39.266747, 39.263355, 39.259968, 39.25658, 39.25319, 39.2498, 39.24921, 39.24862, 39.248028, 39.247437, 39.246845, 39.246254, 39.246834, 39.247414, 39.247993, 39.248573, 39.249153, 39.249733, 39.251995, 39.254257, 39.256523, 39.258785, 39.261047, 39.26331, 39.26784, 39.27237, 39.2769, 39.281433, 39.28596, 39.290493, 39.28993, 39.289368, 39.288803, 39.288242, 39.28768, 39.287117, 39.296185, 39.305256, 39.314323, 39.32339, 39.332462, 39.34153, 39.34436, 39.347195, 39.350025, 39.352856, 39.35569, 39.35852, 39.36644, 39.37436, 39.38228, 39.390198, 39.398117, 39.406036, 39.415115, 39.42419, 39.43327, 39.44235, 39.451424, 39.460503, 39.456528, 39.45255, 39.44857, 39.444595, 39.44062, 39.43664, 39.444584, 39.452526, 39.460472, 39.468414, 39.476357, 39.4843, 39.489975, 39.495647, 39.501324, 39.507, 39.512672, 39.51835, 39.51606, 39.51377, 39.511482, 39.509193, 39.506905, 39.504616, 39.51425, 39.523888, 39.533524, 39.543156, 39.55279, 39.562428, 39.559044, 39.55566, 39.552277, 39.548893, 39.54551, 39.542126, 39.540985, 39.53984, 39.538696, 39.537556, 39.536415, 39.53527, 39.535835, 39.5364, 39.536964, 39.537525, 39.53809, 39.538654, 39.544315, 39.549973, 39.555634, 39.561295, 39.56695, 39.572613, 39.57036, 39.568104, 39.56585, 39.5636, 39.561344, 39.55909, 39.564754, 39.57042, 39.57608, 39.581745, 39.58741, 39.593075, 39.59931, 39.605553, 39.61179, 39.618027, 39.624268, 39.630505, 39.63559, 39.64067, 39.645756, 39.65084, 39.655922, 39.661007, 39.66781, 39.674606, 39.681404, 39.688206, 39.695004, 39.701805, 39.709747, 39.71769, 39.72563, 39.733574, 39.741516, 39.74946, 39.752846, 39.756233, 39.75962, 39.76301, 39.766396, 39.769783, 39.78112, 39.792458, 39.803795, 39.815136, 39.826473, 39.83781, 39.84461, 39.851406, 39.858208, 39.865005, 39.871803, 39.8786, 39.881428, 39.884254, 39.887085, 39.88991, 39.89274, 39.895565, 39.9001, 39.904636, 39.909172, 39.91371, 39.918247, 39.922783, 39.92958, 39.936382, 39.94318, 39.949978, 39.95678, 39.963577, 39.96868, 39.97379, 39.978893, 39.983997, 39.989105, 39.99421, 39.993076, 39.991947, 39.990814, 39.989685, 39.988556, 39.987423, 39.987988, 39.98855, 39.989113, 39.989674, 39.990234, 39.9908, 39.99307, 39.99534, 39.997612, 39.99988, 40.00215, 40.00442, 39.99251, 39.980602, 39.968697, 39.956787, 39.944878, 39.93297, 39.93581, 39.93865, 39.94149, 39.94433, 39.947166, 39.95001, 39.943764, 39.93752, 39.931274, 39.925034, 39.91879, 39.912544, 39.902935, 39.893326, 39.883713, 39.874104, 39.864494, 39.854885, 39.848072, 39.841263, 39.83445, 39.827637, 39.820827, 39.814014, 39.804947, 39.79588, 39.78681, 39.77774, 39.768673, 39.759605, 39.742622, 39.725643, 39.70866, 39.691677, 39.674698, 39.657715, 39.64637, 39.635025, 39.62368, 39.61234, 39.600994, 39.58965, 39.581722, 39.573795, 39.56587, 39.55794, 39.550014, 39.542088, 39.533012, 39.523937, 39.514862, 39.50579, 39.496716, 39.48764, 39.47518, 39.462723, 39.450264, 39.437805, 39.425346, 39.412888, 39.401558, 39.39023, 39.3789, 39.367565, 39.356236, 39.344906, 39.34207, 39.33924, 39.33641, 39.333576, 39.330746, 39.32791, 39.322807, 39.317707, 39.312603, 39.3075, 39.3024, 39.297295, 39.293335, 39.289375, 39.285416, 39.281456, 39.277496, 39.273537, 39.27523, 39.27692, 39.27861, 39.280304, 39.281994, 39.283688, 39.275757, 39.26783, 39.259903, 39.251972, 39.244045, 39.236115, 39.24177, 39.247433, 39.25309, 39.25875, 39.26441, 39.27007, 39.27632, 39.282574, 39.288826, 39.295074, 39.301327, 39.30758, 39.3104, 39.313213, 39.316032, 39.318848, 39.321663, 39.324482, 39.324482, 39.324482, 39.324482, 39.324482, 39.324482, 39.324482, 39.339794, 39.355106, 39.370422, 39.385735, 39.401047, 39.41636, 39.41466, 39.412964, 39.411266, 39.40957, 39.40787, 39.406174, 39.416355, 39.426537, 39.436718, 39.4469, 39.45708, 39.467262, 39.47237, 39.477478, 39.48259, 39.487698, 39.492805, 39.497913, 39.503014, 39.508114, 39.513214, 39.51832, 39.52342, 39.52852, 39.52852, 39.52852, 39.52852, 39.52852, 39.52852, 39.52852, 39.53474, 39.54096, 39.54718, 39.553402, 39.55962, 39.56584, 39.55961, 39.55337, 39.54714, 39.540905, 39.534668, 39.528435, 39.535233, 39.54203, 39.54883, 39.55563, 39.562428, 39.569225, 39.564693, 39.560165, 39.555634, 39.5511, 39.546574, 39.54204, 39.546585, 39.551132, 39.555676, 39.56022, 39.564766, 39.56931, 39.569305, 39.5693, 39.569298, 39.569298, 39.569294, 39.56929, 39.570988, 39.57268, 39.57438, 39.576073, 39.577766, 39.579464, 39.581734, 39.584, 39.58627, 39.58854, 39.590805, 39.593075, 39.600437, 39.607803, 39.615166, 39.62253, 39.629894, 39.63726, 39.642357, 39.64745, 39.652546, 39.657642, 39.662735, 39.66783, 39.67462, 39.68141, 39.6882, 39.694992, 39.701782, 39.708572, 39.71594, 39.72331, 39.730675, 39.738045, 39.74541, 39.75278, 39.74883, 39.744877, 39.74092, 39.73697, 39.733017, 39.729065, 39.744366, 39.759663, 39.774963, 39.790264, 39.80556, 39.82086, 39.830486, 39.840107, 39.84973, 39.859356, 39.868977, 39.8786, 39.8786, 39.8786, 39.8786, 39.8786, 39.8786, 39.8786, 39.887653, 39.89671, 39.90576, 39.914814, 39.92387, 39.932922, 39.93803, 39.943142, 39.94825, 39.953358, 39.95847, 39.963577, 39.965282, 39.966984, 39.96869, 39.97039, 39.97209, 39.973797, 39.97833, 39.982857, 39.98739, 39.991917, 39.996445, 40.000977, 40.00947, 40.01797, 40.026466, 40.03496, 40.04346, 40.051956, 40.047436, 40.042915, 40.038395, 40.033875, 40.029354, 40.024834, 40.01859, 40.01235, 40.006104, 39.999863, 39.99362, 39.987377, 39.981712, 39.976048, 39.970383, 39.964714, 39.95905, 39.953384, 39.948277, 39.943165, 39.938057, 39.93295, 39.927837, 39.92273, 39.917076, 39.911427, 39.905777, 39.900124, 39.894474, 39.88882, 39.876366, 39.86391, 39.851456, 39.839005, 39.82655, 39.814095, 39.80616, 39.79823, 39.7903, 39.782364, 39.774433, 39.7665, 39.756866, 39.747234, 39.737602, 39.727966, 39.718334, 39.708702, 39.6934, 39.678097, 39.662796, 39.647495, 39.63219, 39.61689, 39.61292, 39.60895, 39.60498, 39.601013, 39.597046, 39.593075, 39.5755, 39.55793, 39.54036, 39.522785, 39.505215, 39.48764, 39.478024, 39.468407, 39.45879, 39.449173, 39.439556, 39.42994, 39.42427, 39.418602, 39.412933, 39.40727, 39.4016, 39.39593, 39.387993, 39.380054, 39.372116, 39.364174, 39.356236, 39.348297, 39.344337, 39.340374, 39.33641, 39.33245, 39.32849, 39.324528, 39.326225, 39.327927, 39.329624, 39.33132, 39.333023, 39.33472, 39.325657, 39.316597, 39.307533, 39.298473, 39.289413, 39.28035, 39.28204, 39.28373, 39.28542, 39.28711, 39.2888, 39.29049, 39.28993, 39.289364, 39.288803, 39.288242, 39.287678, 39.287117, 39.289387, 39.291656, 39.293922, 39.296192, 39.298462, 39.30073, 39.303562, 39.306393, 39.309227, 39.312057, 39.314888, 39.31772, 39.327362, 39.337, 39.34664, 39.356285, 39.365925, 39.37557, 39.375553, 39.375538, 39.375523, 39.375507, 39.375492, 39.375477, 39.380013, 39.384552, 39.38909, 39.393627, 39.398163, 39.402702, 39.414597, 39.42649, 39.438385, 39.450283, 39.462177, 39.47407, 39.478615, 39.483154, 39.487698, 39.49224, 39.49678, 39.501324, 39.49622, 39.49111, 39.486008, 39.4809, 39.475796, 39.470688, 39.486546, 39.502407, 39.518265, 39.534122, 39.549984, 39.56584, 39.561874, 39.557907, 39.55394, 39.549976, 39.54601, 39.54204, 39.550537, 39.559036, 39.56753, 39.576027, 39.584526, 39.59302, 39.589634, 39.586246, 39.58286, 39.57947, 39.576084, 39.572697, 39.572697, 39.572697, 39.572697, 39.572697, 39.572697, 39.572697, 39.564754, 39.556816, 39.548874, 39.54093, 39.532993, 39.52505, 39.519955, 39.51486, 39.509758, 39.50466, 39.499565, 39.49447, 39.507504, 39.520535, 39.53357, 39.5466, 39.55963, 39.572666, 39.56756, 39.562447, 39.55734, 39.55223, 39.54712, 39.54201, 39.54995, 39.557888, 39.565826, 39.573765, 39.581703, 39.58964, 39.58681, 39.583984, 39.581154, 39.578323, 39.575497, 39.572666, 39.586273, 39.59988, 39.613487, 39.62709, 39.640697, 39.654305, 39.648632, 39.642956, 39.637283, 39.63161, 39.625935, 39.620262, 39.62706, 39.633858, 39.640656, 39.647457, 39.654255, 39.661053, 39.6656, 39.670147, 39.674698, 39.679245, 39.683792, 39.68834, 39.721752, 39.755165, 39.78858, 39.821995, 39.855408, 39.88882, 39.882595, 39.87637, 39.87014, 39.863914, 39.85769, 39.851463, 39.855415, 39.859367, 39.86332, 39.867268, 39.87122, 39.87517, 39.870087, 39.865, 39.859917, 39.85483, 39.849747, 39.84466, 39.85484, 39.86502, 39.8752, 39.885376, 39.895557, 39.905735, 39.92614, 39.94655, 39.966953, 39.98736, 40.007767, 40.02817, 40.012875, 39.997578, 39.98228, 39.966984, 39.951687, 39.93639, 39.951687, 39.96698, 39.982277, 39.997574, 40.012867, 40.028164, 40.019676, 40.011185, 40.002697, 39.99421, 39.985718, 39.97723, 39.969868, 39.962505, 39.95514, 39.947777, 39.940414, 39.933052, 39.92964, 39.926228, 39.922817, 39.919407, 39.915993, 39.912582, 39.909187, 39.905796, 39.9024, 39.899006, 39.895615, 39.89222, 39.87409, 39.85596, 39.83783, 39.819702, 39.801575, 39.783443, 39.78345, 39.78346, 39.783466, 39.783474, 39.78348, 39.78349, 39.769306, 39.75512, 39.740936, 39.72675, 39.712566, 39.69838, 39.67743, 39.656483, 39.635536, 39.614586, 39.59364, 39.57269, 39.57098, 39.569267, 39.56756, 39.56585, 39.564137, 39.562428, 39.550533, 39.53864, 39.526745, 39.51485, 39.502956, 39.491062, 39.49277, 39.494484, 39.496193, 39.497902, 39.499615, 39.501324, 39.48829, 39.47525, 39.462215, 39.44918, 39.436142, 39.423107, 39.416874, 39.410645, 39.40441, 39.39818, 39.39195, 39.385715, 39.377773, 39.36983, 39.361885, 39.353943, 39.346, 39.33806, 39.336372, 39.33469, 39.333004, 39.331318, 39.329636, 39.32795, 39.333046, 39.338142, 39.34324, 39.348335, 39.35343, 39.35853, 39.361362, 39.364197, 39.367027, 39.36986, 39.372696, 39.37553, 39.369293, 39.363056, 39.35682, 39.35058, 39.34434, 39.338104, 39.328472, 39.31884, 39.309204, 39.299572, 39.28994, 39.280308, 39.292774, 39.30524, 39.317707, 39.330173, 39.34264, 39.355106, 39.353977, 39.35285, 39.351723, 39.350597, 39.349472, 39.348343, 39.34494, 39.341534, 39.33813, 39.33473, 39.33132, 39.32792, 39.33811, 39.34831, 39.3585, 39.368694, 39.37889, 39.389084, 39.39192, 39.39475, 39.397583, 39.400414, 39.403244, 39.40608, 39.422516, 39.438957, 39.4554, 39.471836, 39.488274, 39.504715, 39.503002, 39.50129, 39.499577, 39.497864, 39.49615, 39.49444, 39.49841, 39.50238, 39.50635, 39.510323, 39.514294, 39.518265, 39.51996, 39.521656, 39.52335, 39.525043, 39.52674, 39.528435, 39.526173, 39.523914, 39.521652, 39.51939, 39.51713, 39.51487, 39.519413, 39.523956, 39.528496, 39.53304, 39.537582, 39.542126, 39.54043, 39.538734, 39.537037, 39.53534, 39.533646, 39.531948, 39.5325, 39.533054, 39.533607, 39.534164, 39.534718, 39.53527, 39.530743, 39.52621, 39.521683, 39.517155, 39.512623, 39.508095, 39.507526, 39.506954, 39.506386, 39.505817, 39.505245, 39.504677, 39.50524, 39.505802, 39.506363, 39.506927, 39.50749, 39.508053, 39.51825, 39.528442, 39.53864, 39.548836, 39.55903, 39.569225, 39.56357, 39.557907, 39.552246, 39.54659, 39.54093, 39.53527, 39.538097, 39.540924, 39.543755, 39.54658, 39.549408, 39.552235, 39.559032, 39.56583, 39.572628, 39.579426, 39.586224, 39.59302, 39.60435, 39.615685, 39.627014, 39.638344, 39.649677, 39.661007, 39.667236, 39.673466, 39.679695, 39.68592, 39.69215, 39.69838, 39.712566, 39.72675, 39.740936, 39.75512, 39.769302, 39.78349, 39.78348, 39.783474, 39.783466, 39.78346, 39.78345, 39.783443, 39.784016, 39.784588, 39.785156, 39.78573, 39.7863, 39.786873, 39.7812, 39.77553, 39.76986, 39.76419, 39.758522, 39.75285, 39.763615, 39.77438, 39.785145, 39.79591, 39.806675, 39.81744, 39.824234, 39.831024, 39.83782, 39.844612, 39.851402, 39.858196, 39.850266, 39.842335, 39.834404, 39.826477, 39.818546, 39.810616, 39.819115, 39.82761, 39.83611, 39.84461, 39.853104, 39.861603, 39.855373, 39.849148, 39.84292, 39.836693, 39.830467, 39.824238, 39.81064, 39.79704, 39.78344, 39.76984, 39.75624, 39.74264, 39.75624, 39.76984, 39.78344, 39.79704, 39.81064, 39.824238, 39.819702, 39.815166, 39.81063, 39.806095, 39.80156, 39.797024, 39.783424, 39.769825, 39.756226, 39.742626, 39.729027, 39.715427, 39.705803, 39.69618, 39.686554, 39.676933, 39.66731, 39.657684, 39.657684, 39.65769, 39.65769, 39.65769, 39.657692, 39.657692, 39.654285, 39.650883, 39.647476, 39.64407, 39.640667, 39.63726, 39.631596, 39.625927, 39.620262, 39.614594, 39.60893, 39.60326, 39.58966, 39.57606, 39.56246, 39.548862, 39.535263, 39.521664, 39.509205, 39.496742, 39.484283, 39.471825, 39.459362, 39.446903, 39.439533, 39.43216, 39.42479, 39.417416, 39.410046, 39.40267, 39.414585, 39.4265, 39.438408, 39.45032, 39.462234, 39.474148, 39.456, 39.43786, 39.419712, 39.401566, 39.383423, 39.365276, 39.36415, 39.363026, 39.3619, 39.36078, 39.359653, 39.35853, 39.353428, 39.348324, 39.343224, 39.338123, 39.33302, 39.32792, 39.323387, 39.318855, 39.314323, 39.309795, 39.305264, 39.30073, 39.31092, 39.32111, 39.3313, 39.341484, 39.351673, 39.361862, 39.3545, 39.34714, 39.33978, 39.332417, 39.325058, 39.317696, 39.31599, 39.31428, 39.312576, 39.31087, 39.309162, 39.307457, 39.32446, 39.34146, 39.358463, 39.375465, 39.392467, 39.40947, 39.4191, 39.428734, 39.438366, 39.447998, 39.45763, 39.467262, 39.465572, 39.463882, 39.462196, 39.460506, 39.458817, 39.457127, 39.461655, 39.466183, 39.47071, 39.475243, 39.47977, 39.4843, 39.493366, 39.502434, 39.511505, 39.520573, 39.52964, 39.538708, 39.535313, 39.53192, 39.528526, 39.525135, 39.521744, 39.51835, 39.510983, 39.503616, 39.496246, 39.48888, 39.481514, 39.474148, 39.49114, 39.50813, 39.525116, 39.542107, 39.559097, 39.576088, 39.564747, 39.55341, 39.54207, 39.53073, 39.519394, 39.508053, 39.518257, 39.52846, 39.538666, 39.54887, 39.559074, 39.56928, 39.577213, 39.585148, 39.593086, 39.60102, 39.608955, 39.61689, 39.60386, 39.590828, 39.577797, 39.56477, 39.55174, 39.538708, 39.5336, 39.52849, 39.52338, 39.518272, 39.51316, 39.508053, 39.515423, 39.522797, 39.530167, 39.537537, 39.54491, 39.55228, 39.546036, 39.53979, 39.533546, 39.527306, 39.52106, 39.514816, 39.53183, 39.54884, 39.565853, 39.582867, 39.599876, 39.61689, 39.602726, 39.588562, 39.574394, 39.56023, 39.546066, 39.531902, 39.54096, 39.550014, 39.559074, 39.56813, 39.577187, 39.586243, 39.58002, 39.573795, 39.567574, 39.56135, 39.555126, 39.548904, 39.551174, 39.553444, 39.55571, 39.55798, 39.56025, 39.56252, 39.57611, 39.5897, 39.60329, 39.616882, 39.63047, 39.644062, 39.639534, 39.635006, 39.630478, 39.625946, 39.621418, 39.61689, 39.629345, 39.6418, 39.65426, 39.666714, 39.67917, 39.691624, 39.68652, 39.68142, 39.676315, 39.67121, 39.66611, 39.661007, 39.679714, 39.698418, 39.717125, 39.735832, 39.754536, 39.773243, 39.763607, 39.75397, 39.744335, 39.7347, 39.725063, 39.715427, 39.713165, 39.7109, 39.708637, 39.706375, 39.70411, 39.701847, 39.702984, 39.70412, 39.705254, 39.70639, 39.707527, 39.708664, 39.713764, 39.71887, 39.72397, 39.72907, 39.734173, 39.739273, 39.727924, 39.71658, 39.70523, 39.693886, 39.68254, 39.671192, 39.68027, 39.68935, 39.698425, 39.707504, 39.716583, 39.725662, 39.72962, 39.73358, 39.73754, 39.7415, 39.74546, 39.74942, 39.72959, 39.709763, 39.689934, 39.670105, 39.650276, 39.630447, 39.634407, 39.63837, 39.642334, 39.646294, 39.650253, 39.654217, 39.651947, 39.649677, 39.647408, 39.645138, 39.642868, 39.6406, 39.629276, 39.61795, 39.60663, 39.595306, 39.58398, 39.57266, 39.56417, 39.55568, 39.54719, 39.538704, 39.530212, 39.521725, 39.523983, 39.52624, 39.528496, 39.530754, 39.533012, 39.53527, 39.53131, 39.52735, 39.52339, 39.519436, 39.515476, 39.511517, 39.493942, 39.47637, 39.458797, 39.441223, 39.423653, 39.40608, 39.41061, 39.415142, 39.419678, 39.42421, 39.42874, 39.433273, 39.427048, 39.420826, 39.414604, 39.40838, 39.402157, 39.39593, 39.394234, 39.39254, 39.390842, 39.389145, 39.38745, 39.385754, 39.38404, 39.382328, 39.380615, 39.378902, 39.37719, 39.375477, 39.38059, 39.385696, 39.39081, 39.39592, 39.401028, 39.40614, 39.4016, 39.39706, 39.392517, 39.387978, 39.38344, 39.3789, 39.38626, 39.393623, 39.400986, 39.40835, 39.415714, 39.423077, 39.418545, 39.414013, 39.409485, 39.404953, 39.40042, 39.39589, 39.40213, 39.408367, 39.414608, 39.42085, 39.427086, 39.433327, 39.438427, 39.443527, 39.448624, 39.453724, 39.458824, 39.463924, 39.470158, 39.47639, 39.482624, 39.488857, 39.49509, 39.501324, 39.492825, 39.48432, 39.475822, 39.46732, 39.45882, 39.450317, 39.458813, 39.46731, 39.475807, 39.484303, 39.4928, 39.501297, 39.514896, 39.528496, 39.54209, 39.55569, 39.56929, 39.58289, 39.586857, 39.590824, 39.594788, 39.598755, 39.602722, 39.60669, 39.596478, 39.58627, 39.576057, 39.565845, 39.555637, 39.545425, 39.54317, 39.540916, 39.538666, 39.53641, 39.534157, 39.531902, 39.537567, 39.543232, 39.548897, 39.554558, 39.560223, 39.565887, 39.57042, 39.57495, 39.579483, 39.58401, 39.588543, 39.593075, 39.5857, 39.57833, 39.570957, 39.563583, 39.556213, 39.54884, 39.55338, 39.557922, 39.56246, 39.567005, 39.571545, 39.576088, 39.572124, 39.56816, 39.5642, 39.560238, 39.556274, 39.55231, 39.548904, 39.545494, 39.542088, 39.53868, 39.53527, 39.531864, 39.53527, 39.53868, 39.542088, 39.545494, 39.548904, 39.55231, 39.554012, 39.555714, 39.557415, 39.559116, 39.560818, 39.56252, 39.563644, 39.564774, 39.5659, 39.567024, 39.568153, 39.56928, 39.573246, 39.57721, 39.581177, 39.585144, 39.589108, 39.593075, 39.58628, 39.579487, 39.572693, 39.5659, 39.559105, 39.55231, 39.555702, 39.559097, 39.56249, 39.56588, 39.569275, 39.572666, 39.575512, 39.578354, 39.5812, 39.584045, 39.586887, 39.589733, 39.595966, 39.602196, 39.60843, 39.61466, 39.620888, 39.62712, 39.625977, 39.624836, 39.62369, 39.622547, 39.621407, 39.620262, 39.61912, 39.61798, 39.616844, 39.615704, 39.614563, 39.613422, 39.61627, 39.619118, 39.621964, 39.62481, 39.62766, 39.630505, 39.637867, 39.645226, 39.652588, 39.65995, 39.66731, 39.67467, 39.666733, 39.65879, 39.65085, 39.64291, 39.63497, 39.62703, 39.62137, 39.61571, 39.610054, 39.604393, 39.598736, 39.593075, 39.60158, 39.61009, 39.618595, 39.6271, 39.63561, 39.644115, 39.6356, 39.627083, 39.61857, 39.610054, 39.601536, 39.59302, 39.5868, 39.58058, 39.574364, 39.568142, 39.561924, 39.555702, 39.557972, 39.560238, 39.562508, 39.564774, 39.56704, 39.56931, 39.56647, 39.563633, 39.560795, 39.557957, 39.55512, 39.55228, 39.555668, 39.55906, 39.562447, 39.565834, 39.569225, 39.572613, 39.567524, 39.56244, 39.55735, 39.55226, 39.547176, 39.542088, 39.53813, 39.534176, 39.53022, 39.52626, 39.522305, 39.51835, 39.514942, 39.511536, 39.508133, 39.504726, 39.50132, 39.497913, 39.48375, 39.46959, 39.45543, 39.441265, 39.427105, 39.41294, 39.408974, 39.40501, 39.401043, 39.397076, 39.393112, 39.389145, 39.39934, 39.409534, 39.41973, 39.429928, 39.44012, 39.450317, 39.44296, 39.435604, 39.428246, 39.420887, 39.413532, 39.406174, 39.39937, 39.39256, 39.38575, 39.378944, 39.37214, 39.36533, 39.371555, 39.377777, 39.384003, 39.390224, 39.396446, 39.40267, 39.399273, 39.395878, 39.39248, 39.38908, 39.385685, 39.382286, 39.403816, 39.42535, 39.446884, 39.468414, 39.489944, 39.51148, 39.499004, 39.486534, 39.47406, 39.461586, 39.449116, 39.43664, 39.441196, 39.44575, 39.450306, 39.45486, 39.459415, 39.46397, 39.459423, 39.454876, 39.45033, 39.44578, 39.441235, 39.436687, 39.447456, 39.458225, 39.468994, 39.47976, 39.49053, 39.501297, 39.510357, 39.51942, 39.52848, 39.53754, 39.546604, 39.555664, 39.549995, 39.544327, 39.53866, 39.532993, 39.527325, 39.521656, 39.518826, 39.515995, 39.51317, 39.510338, 39.507507, 39.504677, 39.514317, 39.523956, 39.5336, 39.54324, 39.55288, 39.56252, 39.557972, 39.553425, 39.54888, 39.544334, 39.539787, 39.53524, 39.54771, 39.56018, 39.572655, 39.585125, 39.597595, 39.610065, 39.61063, 39.611195, 39.61176, 39.612324, 39.61289, 39.613453, 39.611763, 39.610077, 39.608387, 39.606697, 39.60501, 39.60332, 39.61011, 39.6169, 39.62369, 39.63048, 39.63727, 39.644062, 39.633865, 39.623672, 39.613476, 39.60328, 39.593086, 39.58289, 39.594215, 39.605545, 39.61687, 39.628197, 39.639526, 39.650852, 39.645752, 39.640656, 39.63556, 39.63046, 39.625362, 39.620262, 39.62196, 39.623657, 39.625355, 39.627052, 39.62875, 39.630447, 39.622517, 39.614582, 39.60665, 39.598717, 39.590786, 39.58285, 39.581154, 39.579456, 39.57776, 39.57606, 39.574364, 39.572666, 39.580044, 39.58742, 39.594795, 39.602173, 39.60955, 39.61693, 39.62598, 39.635033, 39.64408, 39.653133, 39.662186, 39.671238, 39.666138, 39.66104, 39.655945, 39.650845, 39.64575, 39.640648, 39.635544, 39.63044, 39.625336, 39.620235, 39.61513, 39.610027, 39.607193, 39.60436, 39.601524, 39.59869, 39.595856, 39.59302, 39.597008, 39.60099, 39.604973, 39.60896, 39.61294, 39.61693, 39.615223, 39.613514, 39.61181, 39.610104, 39.608395, 39.60669, 39.606117, 39.605545, 39.604973, 39.604404, 39.603832, 39.60326, 39.59307, 39.582882, 39.572693, 39.562504, 39.552315, 39.542126, 39.55006, 39.557995, 39.56593, 39.573864, 39.5818, 39.589733, 39.572155, 39.554573, 39.536995, 39.519413, 39.501835, 39.484253, 39.497284, 39.51031, 39.52334, 39.53637, 39.549397, 39.562428, 39.551666, 39.54091, 39.530148, 39.519386, 39.50863, 39.497868, 39.504665, 39.511463, 39.51826, 39.52506, 39.531857, 39.538654, 39.537514, 39.536373, 39.535233, 39.534092, 39.53295, 39.53181, 39.525585, 39.519363, 39.513138, 39.506916, 39.500694, 39.49447, 39.49673, 39.498997, 39.50126, 39.503525, 39.505787, 39.508053, 39.50748, 39.50691, 39.506332, 39.50576, 39.505188, 39.504616, 39.49727, 39.489925, 39.48258, 39.47523, 39.467888, 39.46054, 39.461662, 39.46278, 39.4639, 39.465023, 39.46614, 39.467262, 39.459343, 39.451427, 39.44351, 39.43559, 39.427673, 39.419754, 39.41578, 39.411804, 39.40783, 39.40385, 39.399876, 39.3959, 39.392498, 39.38909, 39.38569, 39.382286, 39.37888, 39.375477, 39.38115, 39.38682, 39.392494, 39.39817, 39.403843, 39.409515, 39.40555, 39.401577, 39.39761, 39.393642, 39.38967, 39.385704, 39.389107, 39.392513, 39.39592, 39.399323, 39.402725, 39.40613, 39.402725, 39.399323, 39.39592, 39.392513, 39.38911, 39.385704, 39.389114, 39.39253, 39.39594, 39.39935, 39.402763, 39.406174, 39.40956, 39.41295, 39.416336, 39.419727, 39.423115, 39.426502, 39.42933, 39.432156, 39.434982, 39.43781, 39.440636, 39.443462, 39.45367, 39.46388, 39.47409, 39.4843, 39.494507, 39.504715, 39.499603, 39.494488, 39.489372, 39.48426, 39.47915, 39.474033, 39.480274, 39.486515, 39.492756, 39.498997, 39.505238, 39.51148, 39.517136, 39.522793, 39.52845, 39.53411, 39.53977, 39.545425, 39.548264, 39.5511, 39.55394, 39.556778, 39.559616, 39.562454, 39.561893, 39.561333, 39.560772, 39.56021, 39.55965, 39.55909, 39.56078, 39.56247, 39.564156, 39.565845, 39.567535, 39.569225, 39.57036, 39.57149, 39.572624, 39.57376, 39.574894, 39.576027, 39.58227, 39.588516, 39.594757, 39.601, 39.607246, 39.61349, 39.61462, 39.61575, 39.616875, 39.618004, 39.619133, 39.620262, 39.621967, 39.623676, 39.62538, 39.627087, 39.628796, 39.6305, 39.629356, 39.628216, 39.627075, 39.62593, 39.62479, 39.623646, 39.62479, 39.62593, 39.627075, 39.62822, 39.62936, 39.630505, 39.629368, 39.62823, 39.62709, 39.625954, 39.624817, 39.62368, 39.624817, 39.625954, 39.62709, 39.628227, 39.629364, 39.6305, 39.62992, 39.629345, 39.628765, 39.628185, 39.62761, 39.62703, 39.631, 39.63497, 39.638947, 39.642918, 39.64689, 39.65086, 39.645203, 39.63955, 39.633896, 39.62824, 39.622585, 39.61693, 39.615223, 39.613514, 39.61181, 39.610104, 39.608395, 39.60669, 39.610664, 39.614635, 39.61861, 39.622585, 39.626556, 39.63053, 39.630527, 39.630524, 39.630516, 39.630512, 39.63051, 39.630505, 39.627098, 39.62369, 39.620285, 39.61688, 39.613472, 39.610065, 39.608364, 39.60666, 39.604958, 39.603252, 39.60155, 39.599846, 39.600418, 39.600986, 39.601555, 39.602127, 39.602695, 39.603268, 39.601013, 39.598755, 39.5965, 39.594246, 39.591988, 39.589733, 39.588593, 39.587452, 39.58631, 39.58517, 39.58403, 39.58289, 39.57666, 39.57043, 39.5642, 39.55797, 39.55174, 39.54551, 39.5421, 39.53869, 39.53528, 39.53187, 39.52846, 39.52505, 39.521656, 39.51826, 39.514862, 39.511467, 39.50807, 39.504677, 39.499588, 39.4945, 39.48941, 39.484325, 39.479237, 39.474148, 39.474148, 39.474148, 39.474148, 39.474148, 39.474148, 39.474148, 39.473007, 39.471863, 39.470722, 39.46958, 39.468437, 39.467297, 39.460506, 39.453716, 39.446926, 39.440136, 39.433346, 39.426556, 39.42258, 39.418606, 39.414627, 39.410652, 39.406677, 39.402702, 39.398727, 39.394753, 39.390778, 39.386803, 39.382828, 39.378853, 39.376606, 39.37436, 39.372116, 39.36987, 39.367622, 39.365376, 39.368195, 39.371014, 39.373833, 39.376648, 39.379467, 39.382286, 39.37662, 39.370956, 39.36529, 39.359627, 39.353962, 39.348297, 39.347164, 39.34603, 39.344894, 39.34376, 39.34263, 39.341496, 39.34093, 39.340366, 39.339798, 39.339233, 39.33867, 39.338104, 39.338104, 39.338104, 39.338104, 39.338104, 39.338104, 39.338104, 39.338097, 39.33809, 39.33808, 39.338074, 39.338066, 39.33806, 39.33977, 39.341488, 39.3432, 39.344913, 39.34663, 39.348343, 39.351738, 39.355133, 39.35853, 39.361923, 39.36532, 39.368713, 39.367584, 39.36646, 39.365334, 39.364204, 39.36308, 39.36195, 39.364204, 39.36646, 39.368713, 39.370968, 39.373222, 39.375477, 39.37888, 39.382282, 39.38568, 39.389084, 39.392487, 39.39589, 39.39985, 39.403812, 39.407772, 39.41173, 39.415695, 39.419655, 39.425888, 39.432117, 39.438347, 39.44458, 39.45081, 39.457043, 39.459873, 39.462708, 39.465538, 39.46837, 39.471203, 39.474033, 39.478577, 39.48312, 39.487663, 39.492207, 39.49675, 39.501293, 39.50638, 39.511467, 39.516552, 39.521637, 39.526726, 39.53181, 39.528988, 39.526165, 39.52334, 39.520515, 39.517693, 39.51487, 39.521675, 39.52848, 39.535286, 39.54209, 39.548897, 39.555702, 39.555687, 39.555676, 39.555664, 39.55565, 39.555637, 39.555622, 39.56356, 39.571503, 39.57944, 39.58738, 39.59532, 39.60326, 39.598167, 39.59307, 39.58798, 39.582886, 39.57779, 39.572697, 39.57609, 39.57949, 39.582886, 39.58628, 39.58968, 39.593075, 39.59705, 39.601025, 39.605003, 39.60898, 39.612953, 39.61693, 39.614082, 39.611233, 39.608387, 39.60554, 39.60269, 39.599846, 39.60721, 39.614567, 39.621925, 39.629288, 39.636646, 39.64401, 39.64911, 39.654213, 39.659313, 39.664413, 39.669518, 39.674618, 39.676907, 39.67919, 39.68148, 39.683765, 39.68605, 39.68834, 39.683784, 39.67923, 39.674675, 39.670116, 39.66556, 39.661007, 39.667812, 39.67462, 39.681427, 39.688232, 39.69504, 39.701847, 39.69957, 39.697296, 39.695023, 39.692745, 39.69047, 39.688194, 39.683098, 39.678005, 39.67291, 39.667812, 39.66272, 39.657623, 39.658188, 39.658752, 39.659317, 39.659878, 39.660442, 39.661007, 39.658752, 39.656498, 39.654243, 39.651993, 39.64974, 39.647484, 39.647484, 39.647484, 39.647484, 39.647484, 39.647484, 39.647484, 39.645786, 39.644085, 39.642387, 39.64069, 39.63899, 39.63729, 39.634457, 39.631622, 39.62879, 39.625957, 39.623123, 39.62029, 39.618584, 39.616882, 39.615177, 39.613472, 39.61177, 39.610065, 39.609493, 39.60892, 39.608353, 39.60778, 39.60721, 39.606636, 39.59814, 39.589645, 39.58115, 39.572655, 39.56416, 39.555664, 39.55454, 39.55341, 39.552284, 39.55116, 39.55003, 39.548904, 39.543224, 39.53754, 39.53186, 39.52618, 39.520496, 39.514816, 39.517673, 39.520527, 39.523384, 39.526237, 39.52909, 39.531948, 39.524563, 39.517178, 39.509796, 39.50241, 39.495026, 39.48764, 39.478024, 39.468407, 39.45879, 39.449173, 39.439556, 39.42994, 39.42313, 39.416325, 39.409515, 39.402706, 39.3959, 39.38909, 39.389088, 39.38908, 39.389076, 39.389072, 39.389065, 39.38906, 39.383957, 39.378853, 39.37375, 39.368645, 39.36354, 39.358437, 39.356747, 39.355057, 39.353367, 39.351677, 39.349987, 39.348297, 39.348858, 39.34942, 39.349983, 39.350544, 39.351105, 39.351665, 39.346004, 39.34034, 39.33468, 39.329014, 39.323353, 39.317688, 39.317688, 39.31769, 39.31769, 39.31769, 39.317696, 39.317696, 39.3126, 39.307503, 39.302406, 39.29731, 39.292213, 39.287117, 39.287678, 39.288242, 39.288803, 39.289364, 39.28993, 39.29049, 39.297863, 39.305233, 39.312607, 39.319977, 39.327347, 39.33472, 39.335278, 39.335835, 39.336388, 39.336945, 39.3375, 39.33806, 39.344303, 39.35055, 39.356796, 39.36304, 39.36929, 39.375534, 39.378925, 39.38232, 39.38571, 39.389103, 39.392498, 39.39589, 39.3993, 39.402714, 39.406124, 39.409534, 39.41295, 39.41636, 39.42258, 39.428802, 39.43502, 39.441242, 39.447464, 39.453686, 39.457092, 39.460495, 39.4639, 39.467308, 39.47071, 39.474117, 39.47412, 39.47413, 39.474133, 39.474136, 39.474144, 39.474148, 39.483196, 39.492245, 39.50129, 39.510338, 39.519386, 39.528435, 39.530712, 39.532986, 39.535263, 39.537537, 39.53981, 39.542088, 39.545483, 39.548874, 39.55227, 39.555664, 39.559055, 39.56245, 39.56812, 39.573788, 39.57946, 39.58513, 39.590797, 39.596466, 38.02403, 36.45159, 34.879158, 33.30672, 31.734283, 30.161848, 24.922405, 19.682962, 14.44352, 9.204076, 3.964634, -1.2748094, -1.2759597, -1.27711, -1.2782602, -1.2794106, -1.280561, -1.2817112, -1.2828573, -1.2840033, -1.2851493, -1.2862954, -1.2874415, -1.2885876, -1.2908757, -1.2931638, -1.2954519, -1.29774, -1.3000281, -1.3023162, -1.3063213, -1.3103263, -1.3143315, -1.3183365, -1.3223417, -1.3263468, -1.3269219, -1.327497, -1.3280722, -1.3286474, -1.3292226, -1.3297977, -1.3320868, -1.3343759, -1.3366649, -1.338954}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
