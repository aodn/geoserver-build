netcdf file-129.nc {
  dimensions:
    DEPTH = 29;
  variables:
    float LATITUDE(DEPTH=29);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=29);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=29);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=29);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=29);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=29);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593, 23061.036030092593}
TEMP =
  {28.8775, 28.7094, 28.6336, 28.5961, 28.5701, 28.5469, 28.5256, 28.5093, 28.5045, 28.4978, 28.4907, 28.4767, 28.4667, 28.4606, 28.4584, 28.4597, 28.4545, 28.4525, 28.4512, 28.4499, 28.4503, 28.4486, 28.4491, 28.4494, 28.4494, 28.4492, 28.4504, 28.4535, 28.4555}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829, 28.823}
}
