netcdf file-168.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (29 currently)
  variables:
    float LATITUDE(DEPTH=29);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=29);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=29);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=29);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=29);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=29);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962, 22656.086400462962}
TEMP =
  {28.8875, 28.8085, 28.776, 28.7894, 28.7746, 28.7481, 28.7116, 28.7021, 28.7096, 28.6834, 28.663, 28.6583, 28.659, 28.6553, 28.6532, 28.6519, 28.6505, 28.6509, 28.6508, 28.6495, 28.6486, 28.6488, 28.649, 28.6483, 28.6481, 28.6482, 28.6487, 28.649, 28.6492}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829, 28.823}
}
