netcdf file-162.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (17 currently)
  variables:
    float LATITUDE(DEPTH=17);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=17);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=17);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=17);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=17);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=17);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296, 22446.034733796296}
TEMP =
  {22.6664, 22.665, 22.6638, 22.6629, 22.6623, 22.662, 22.6616, 22.661, 22.6608, 22.6606, 22.6606, 22.661, 22.6608, 22.6602, 22.6599, 22.66, 22.6603}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.902, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853}
}
