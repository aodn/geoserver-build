netcdf file-159.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (23 currently)
  variables:
    float LATITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=23);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=23);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=23);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=23);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926, 22361.045613425926}
TEMP =
  {28.6137, 28.5154, 28.4375, 28.387, 28.346, 28.3013, 28.2474, 28.1849, 28.1203, 28.0539, 27.9771, 27.8986, 27.8302, 27.7694, 27.7136, 27.6769, 27.6553, 27.64, 27.6308, 27.6263, 27.6245, 27.624, 27.6236}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.982, 3.976, 4.969, 5.964, 6.958, 7.951, 8.946, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847}
}
