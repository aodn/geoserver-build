netcdf file-171.nc {
  dimensions:
    DEPTH = 28;
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193, 147.6193}
TIME =
  {22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185, 22759.046747685185}
TEMP =
  {26.8903, 26.8654, 26.8489, 26.8303, 26.8133, 26.8027, 26.7968, 26.7947, 26.7945, 26.7942, 26.7929, 26.7903, 26.7894, 26.789, 26.7898, 26.7923, 26.7946, 26.7967, 26.8016, 26.8122, 26.8246, 26.8288, 26.83, 26.8318, 26.8332, 26.834, 26.8349, 26.8351}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
