netcdf file-116.nc {
  dimensions:
    DEPTH = 20;
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297, 22987.895046296297}
TEMP =
  {31.8905, 31.8922, 31.8928, 31.8959, 31.8973, 31.8973, 31.8975, 31.8977, 31.8977, 31.898, 31.8984, 31.8981, 31.8984, 31.8993, 31.8996, 31.8998, 31.8998, 31.9008, 31.9031, 31.9031}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879}
}
