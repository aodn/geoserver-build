netcdf file-47.nc {
  dimensions:
    DEPTH = 43;
  variables:
    float LATITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=43);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=43);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223, 22674.156597222223}
TEMP =
  {23.5187, 23.5212, 23.5189, 23.5176, 23.5158, 23.5117, 23.5104, 23.5112, 23.5095, 23.508, 23.5067, 23.5039, 23.5061, 23.5115, 23.5198, 23.5204, 23.5193, 23.517, 23.5056, 23.4988, 23.4978, 23.4915, 23.4886, 23.4817, 23.4713, 23.4585, 23.4349, 23.2944, 23.069, 22.6538, 22.2077, 22.1068, 22.0395, 22.0085, 21.9822, 21.9707, 21.9607, 21.9544, 21.9583, 21.9334, 21.9153, 21.906, 21.9022}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0}
}
