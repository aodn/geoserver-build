netcdf file-161.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (24 currently)
  variables:
    float LATITUDE(DEPTH=24);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=24);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=24);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=24);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=24);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=24);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705, 22426.040266203705}
TEMP =
  {23.5981, 23.6012, 23.6044, 23.6078, 23.6082, 23.6086, 23.6092, 23.6093, 23.609, 23.6083, 23.6085, 23.6082, 23.609, 23.6096, 23.6103, 23.6107, 23.6109, 23.6104, 23.6096, 23.6093, 23.6094, 23.6094, 23.6094, 23.6099}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853}
}
