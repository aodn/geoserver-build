netcdf file-92.nc {
  dimensions:
    DEPTH = 21;
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556, 23178.771805555556}
TEMP =
  {26.9847, 26.9872, 26.9871, 26.9865, 26.9868, 26.9888, 26.9884, 26.9879, 26.9881, 26.9885, 26.9774, 26.9809, 26.9795, 26.9835, 26.9881, 26.9899, 26.9905, 26.9905, 26.9906, 26.9907, 26.9891}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872}
}
