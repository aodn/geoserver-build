netcdf IMOS_ANMN-TS_20150113T230000Z_WATR20_FV01_WATR20-1407-Nortek-ADCP-190kHz-194_END-20150121T021500Z_id-7736.nc {
  dimensions:
    TIME = UNLIMITED;   // (686 currently)
  variables:
    double TIME(TIME=686);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=686);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=686);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=686);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=686);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=686);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=686);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=686);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=686);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=686);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=686);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=686);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=686);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical max information has been computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :instrument = "Nortek       ADCP 190kHz";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "CNL6105";
  :history = "2015-01-29T06:31:59Z - depthPP: Depth computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).\n2015-01-29T06:32:03Z - magneticDeclinationPP: data initially referring to magnetic North has been modified so that it now refers to true North, applying a computed magnetic declination of -1.9667degrees. NOAA\'s Geomag v7.0 software + IGRF11 model have been used to compute this value at a latitude=-31.7286degrees North, longitude=115.0371degrees East, depth=194m (instrument nominal depth) and date=2014/10/15 (date in the middle of time_coverage_start and time_coverage_end).";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 194.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = 0.3984445f; // float
  :geospatial_vertical_max = 206.16779f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-21T02:15:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.96875, 23753.979166666668, 23753.989583333332, 23754.0, 23754.010416666668, 23754.020833333332, 23754.03125, 23754.041666666668, 23754.052083333332, 23754.0625, 23754.072916666668, 23754.083333333332, 23754.09375, 23754.104166666668, 23754.114583333332, 23754.125, 23754.135416666668, 23754.145833333332, 23754.15625, 23754.166666666668, 23754.177083333332, 23754.1875, 23754.197916666668, 23754.208333333332, 23754.21875, 23754.229166666668, 23754.239583333332, 23754.25, 23754.260416666668, 23754.270833333332, 23754.28125, 23754.291666666668, 23754.302083333332, 23754.3125, 23754.322916666668, 23754.333333333332, 23754.34375, 23754.354166666668, 23754.364583333332, 23754.375, 23754.385416666668, 23754.395833333332, 23754.40625, 23754.416666666668, 23754.427083333332, 23754.4375, 23754.447916666668, 23754.458333333332, 23754.46875, 23754.479166666668, 23754.489583333332, 23754.5, 23754.510416666668, 23754.520833333332, 23754.53125, 23754.541666666668, 23754.552083333332, 23754.5625, 23754.572916666668, 23754.583333333332, 23754.59375, 23754.604166666668, 23754.614583333332, 23754.625, 23754.635416666668, 23754.645833333332, 23754.65625, 23754.666666666668, 23754.677083333332, 23754.6875, 23754.697916666668, 23754.708333333332, 23754.71875, 23754.729166666668, 23754.739583333332, 23754.75, 23754.760416666668, 23754.770833333332, 23754.78125, 23754.791666666668, 23754.802083333332, 23754.8125, 23754.822916666668, 23754.833333333332, 23754.84375, 23754.854166666668, 23754.864583333332, 23754.875, 23754.885416666668, 23754.895833333332, 23754.90625, 23754.916666666668, 23754.927083333332, 23754.9375, 23754.947916666668, 23754.958333333332, 23754.96875, 23754.979166666668, 23754.989583333332, 23755.0, 23755.010416666668, 23755.020833333332, 23755.03125, 23755.041666666668, 23755.052083333332, 23755.0625, 23755.072916666668, 23755.083333333332, 23755.09375, 23755.104166666668, 23755.114583333332, 23755.125, 23755.135416666668, 23755.145833333332, 23755.15625, 23755.166666666668, 23755.177083333332, 23755.1875, 23755.197916666668, 23755.208333333332, 23755.21875, 23755.229166666668, 23755.239583333332, 23755.25, 23755.260416666668, 23755.270833333332, 23755.28125, 23755.291666666668, 23755.302083333332, 23755.3125, 23755.322916666668, 23755.333333333332, 23755.34375, 23755.354166666668, 23755.364583333332, 23755.375, 23755.385416666668, 23755.395833333332, 23755.40625, 23755.416666666668, 23755.427083333332, 23755.4375, 23755.447916666668, 23755.458333333332, 23755.46875, 23755.479166666668, 23755.489583333332, 23755.5, 23755.510416666668, 23755.520833333332, 23755.53125, 23755.541666666668, 23755.552083333332, 23755.5625, 23755.572916666668, 23755.583333333332, 23755.59375, 23755.604166666668, 23755.614583333332, 23755.625, 23755.635416666668, 23755.645833333332, 23755.65625, 23755.666666666668, 23755.677083333332, 23755.6875, 23755.697916666668, 23755.708333333332, 23755.71875, 23755.729166666668, 23755.739583333332, 23755.75, 23755.760416666668, 23755.770833333332, 23755.78125, 23755.791666666668, 23755.802083333332, 23755.8125, 23755.822916666668, 23755.833333333332, 23755.84375, 23755.854166666668, 23755.864583333332, 23755.875, 23755.885416666668, 23755.895833333332, 23755.90625, 23755.916666666668, 23755.927083333332, 23755.9375, 23755.947916666668, 23755.958333333332, 23755.96875, 23755.979166666668, 23755.989583333332, 23756.0, 23756.010416666668, 23756.020833333332, 23756.03125, 23756.041666666668, 23756.052083333332, 23756.0625, 23756.072916666668, 23756.083333333332, 23756.09375, 23756.104166666668, 23756.114583333332, 23756.125, 23756.135416666668, 23756.145833333332, 23756.15625, 23756.166666666668, 23756.177083333332, 23756.1875, 23756.197916666668, 23756.208333333332, 23756.21875, 23756.229166666668, 23756.239583333332, 23756.25, 23756.260416666668, 23756.270833333332, 23756.28125, 23756.291666666668, 23756.302083333332, 23756.3125, 23756.322916666668, 23756.333333333332, 23756.34375, 23756.354166666668, 23756.364583333332, 23756.375, 23756.385416666668, 23756.395833333332, 23756.40625, 23756.416666666668, 23756.427083333332, 23756.4375, 23756.447916666668, 23756.458333333332, 23756.46875, 23756.479166666668, 23756.489583333332, 23756.5, 23756.510416666668, 23756.520833333332, 23756.53125, 23756.541666666668, 23756.552083333332, 23756.5625, 23756.572916666668, 23756.583333333332, 23756.59375, 23756.604166666668, 23756.614583333332, 23756.625, 23756.635416666668, 23756.645833333332, 23756.65625, 23756.666666666668, 23756.677083333332, 23756.6875, 23756.697916666668, 23756.708333333332, 23756.71875, 23756.729166666668, 23756.739583333332, 23756.75, 23756.760416666668, 23756.770833333332, 23756.78125, 23756.791666666668, 23756.802083333332, 23756.8125, 23756.822916666668, 23756.833333333332, 23756.84375, 23756.854166666668, 23756.864583333332, 23756.875, 23756.885416666668, 23756.895833333332, 23756.90625, 23756.916666666668, 23756.927083333332, 23756.9375, 23756.947916666668, 23756.958333333332, 23756.96875, 23756.979166666668, 23756.989583333332, 23757.0, 23757.010416666668, 23757.020833333332, 23757.03125, 23757.041666666668, 23757.052083333332, 23757.0625, 23757.072916666668, 23757.083333333332, 23757.09375, 23757.104166666668, 23757.114583333332, 23757.125, 23757.135416666668, 23757.145833333332, 23757.15625, 23757.166666666668, 23757.177083333332, 23757.1875, 23757.197916666668, 23757.208333333332, 23757.21875, 23757.229166666668, 23757.239583333332, 23757.25, 23757.260416666668, 23757.270833333332, 23757.28125, 23757.291666666668, 23757.302083333332, 23757.3125, 23757.322916666668, 23757.333333333332, 23757.34375, 23757.354166666668, 23757.364583333332, 23757.375, 23757.385416666668, 23757.395833333332, 23757.40625, 23757.416666666668, 23757.427083333332, 23757.4375, 23757.447916666668, 23757.458333333332, 23757.46875, 23757.479166666668, 23757.489583333332, 23757.5, 23757.510416666668, 23757.520833333332, 23757.53125, 23757.541666666668, 23757.552083333332, 23757.5625, 23757.572916666668, 23757.583333333332, 23757.59375, 23757.604166666668, 23757.614583333332, 23757.625, 23757.635416666668, 23757.645833333332, 23757.65625, 23757.666666666668, 23757.677083333332, 23757.6875, 23757.697916666668, 23757.708333333332, 23757.71875, 23757.729166666668, 23757.739583333332, 23757.75, 23757.760416666668, 23757.770833333332, 23757.78125, 23757.791666666668, 23757.802083333332, 23757.8125, 23757.822916666668, 23757.833333333332, 23757.84375, 23757.854166666668, 23757.864583333332, 23757.875, 23757.885416666668, 23757.895833333332, 23757.90625, 23757.916666666668, 23757.927083333332, 23757.9375, 23757.947916666668, 23757.958333333332, 23757.96875, 23757.979166666668, 23757.989583333332, 23758.0, 23758.010416666668, 23758.020833333332, 23758.03125, 23758.041666666668, 23758.052083333332, 23758.0625, 23758.072916666668, 23758.083333333332, 23758.09375, 23758.104166666668, 23758.114583333332, 23758.125, 23758.135416666668, 23758.145833333332, 23758.15625, 23758.166666666668, 23758.177083333332, 23758.1875, 23758.197916666668, 23758.208333333332, 23758.21875, 23758.229166666668, 23758.239583333332, 23758.25, 23758.260416666668, 23758.270833333332, 23758.28125, 23758.291666666668, 23758.302083333332, 23758.3125, 23758.322916666668, 23758.333333333332, 23758.34375, 23758.354166666668, 23758.364583333332, 23758.375, 23758.385416666668, 23758.395833333332, 23758.40625, 23758.416666666668, 23758.427083333332, 23758.4375, 23758.447916666668, 23758.458333333332, 23758.46875, 23758.479166666668, 23758.489583333332, 23758.5, 23758.510416666668, 23758.520833333332, 23758.53125, 23758.541666666668, 23758.552083333332, 23758.5625, 23758.572916666668, 23758.583333333332, 23758.59375, 23758.604166666668, 23758.614583333332, 23758.625, 23758.635416666668, 23758.645833333332, 23758.65625, 23758.666666666668, 23758.677083333332, 23758.6875, 23758.697916666668, 23758.708333333332, 23758.71875, 23758.729166666668, 23758.739583333332, 23758.75, 23758.760416666668, 23758.770833333332, 23758.78125, 23758.791666666668, 23758.802083333332, 23758.8125, 23758.822916666668, 23758.833333333332, 23758.84375, 23758.854166666668, 23758.864583333332, 23758.875, 23758.885416666668, 23758.895833333332, 23758.90625, 23758.916666666668, 23758.927083333332, 23758.9375, 23758.947916666668, 23758.958333333332, 23758.96875, 23758.979166666668, 23758.989583333332, 23759.0, 23759.010416666668, 23759.020833333332, 23759.03125, 23759.041666666668, 23759.052083333332, 23759.0625, 23759.072916666668, 23759.083333333332, 23759.09375, 23759.104166666668, 23759.114583333332, 23759.125, 23759.135416666668, 23759.145833333332, 23759.15625, 23759.166666666668, 23759.177083333332, 23759.1875, 23759.197916666668, 23759.208333333332, 23759.21875, 23759.229166666668, 23759.239583333332, 23759.25, 23759.260416666668, 23759.270833333332, 23759.28125, 23759.291666666668, 23759.302083333332, 23759.3125, 23759.322916666668, 23759.333333333332, 23759.34375, 23759.354166666668, 23759.364583333332, 23759.375, 23759.385416666668, 23759.395833333332, 23759.40625, 23759.416666666668, 23759.427083333332, 23759.4375, 23759.447916666668, 23759.458333333332, 23759.46875, 23759.479166666668, 23759.489583333332, 23759.5, 23759.510416666668, 23759.520833333332, 23759.53125, 23759.541666666668, 23759.552083333332, 23759.5625, 23759.572916666668, 23759.583333333332, 23759.59375, 23759.604166666668, 23759.614583333332, 23759.625, 23759.635416666668, 23759.645833333332, 23759.65625, 23759.666666666668, 23759.677083333332, 23759.6875, 23759.697916666668, 23759.708333333332, 23759.71875, 23759.729166666668, 23759.739583333332, 23759.75, 23759.760416666668, 23759.770833333332, 23759.78125, 23759.791666666668, 23759.802083333332, 23759.8125, 23759.822916666668, 23759.833333333332, 23759.84375, 23759.854166666668, 23759.864583333332, 23759.875, 23759.885416666668, 23759.895833333332, 23759.90625, 23759.916666666668, 23759.927083333332, 23759.9375, 23759.947916666668, 23759.958333333332, 23759.96875, 23759.979166666668, 23759.989583333332, 23760.0, 23760.010416666668, 23760.020833333332, 23760.03125, 23760.041666666668, 23760.052083333332, 23760.0625, 23760.072916666668, 23760.083333333332, 23760.09375, 23760.104166666668, 23760.114583333332, 23760.125, 23760.135416666668, 23760.145833333332, 23760.15625, 23760.166666666668, 23760.177083333332, 23760.1875, 23760.197916666668, 23760.208333333332, 23760.21875, 23760.229166666668, 23760.239583333332, 23760.25, 23760.260416666668, 23760.270833333332, 23760.28125, 23760.291666666668, 23760.302083333332, 23760.3125, 23760.322916666668, 23760.333333333332, 23760.34375, 23760.354166666668, 23760.364583333332, 23760.375, 23760.385416666668, 23760.395833333332, 23760.40625, 23760.416666666668, 23760.427083333332, 23760.4375, 23760.447916666668, 23760.458333333332, 23760.46875, 23760.479166666668, 23760.489583333332, 23760.5, 23760.510416666668, 23760.520833333332, 23760.53125, 23760.541666666668, 23760.552083333332, 23760.5625, 23760.572916666668, 23760.583333333332, 23760.59375, 23760.604166666668, 23760.614583333332, 23760.625, 23760.635416666668, 23760.645833333332, 23760.65625, 23760.666666666668, 23760.677083333332, 23760.6875, 23760.697916666668, 23760.708333333332, 23760.71875, 23760.729166666668, 23760.739583333332, 23760.75, 23760.760416666668, 23760.770833333332, 23760.78125, 23760.791666666668, 23760.802083333332, 23760.8125, 23760.822916666668, 23760.833333333332, 23760.84375, 23760.854166666668, 23760.864583333332, 23760.875, 23760.885416666668, 23760.895833333332, 23760.90625, 23760.916666666668, 23760.927083333332, 23760.9375, 23760.947916666668, 23760.958333333332, 23760.96875, 23760.979166666668, 23760.989583333332, 23761.0, 23761.010416666668, 23761.020833333332, 23761.03125, 23761.041666666668, 23761.052083333332, 23761.0625, 23761.072916666668, 23761.083333333332, 23761.09375}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =194.0
TEMP =
  {16.33, 16.29, 16.24, 16.19, 16.14, 16.1, 16.07, 16.03, 15.99, 15.95, 15.92, 15.89, 15.88, 15.89, 15.92, 15.98, 16.05, 16.14, 16.22, 16.29, 16.35, 16.4, 16.43, 16.45, 16.47, 16.48, 16.5, 16.51, 16.52, 16.53, 16.55, 16.57, 16.59, 16.61, 16.63, 16.64, 16.66, 16.67, 16.69, 16.7, 16.71, 16.71, 16.72, 16.72, 16.72, 16.72, 16.71, 16.7, 16.7, 16.7, 16.7, 16.71, 16.71, 16.72, 16.72, 16.74, 16.74, 16.75, 16.75, 16.76, 16.76, 16.77, 16.78, 16.79, 16.8, 16.81, 16.82, 16.83, 16.85, 16.86, 16.87, 16.88, 16.88, 16.89, 16.9, 16.91, 16.93, 16.94, 16.96, 16.97, 16.99, 17.01, 17.03, 17.06, 17.09, 17.11, 17.14, 17.16, 17.17, 17.19, 17.17, 17.08, 16.94, 16.73, 16.51, 16.29, 16.11, 15.95, 15.82, 15.72, 15.63, 15.56, 15.5, 15.45, 15.44, 15.48, 15.56, 15.69, 15.86, 16.04, 16.21, 16.37, 16.51, 16.62, 16.71, 16.78, 16.81, 16.82, 16.83, 16.85, 16.88, 16.91, 16.96, 17.01, 17.07, 17.13, 17.18, 17.22, 17.26, 17.3, 17.33, 17.35, 17.37, 17.38, 17.39, 17.39, 17.4, 17.41, 17.42, 17.43, 17.44, 17.45, 17.46, 17.45, 17.45, 17.45, 17.45, 17.45, 17.46, 17.44, 17.39, 17.34, 17.3, 17.27, 17.24, 17.21, 17.19, 17.18, 17.19, 17.21, 17.24, 17.27, 17.28, 17.3, 17.32, 17.32, 17.34, 17.35, 17.37, 17.39, 17.41, 17.42, 17.44, 17.46, 17.48, 17.5, 17.52, 17.54, 17.56, 17.58, 17.59, 17.57, 17.46, 17.23, 16.85, 16.38, 15.92, 15.54, 15.21, 14.94, 14.72, 14.55, 14.42, 14.31, 14.21, 14.12, 14.04, 13.97, 13.91, 13.86, 13.82, 13.79, 13.78, 13.79, 13.81, 13.85, 13.89, 13.93, 13.97, 14.03, 14.13, 14.28, 14.49, 14.72, 14.94, 15.21, 15.53, 15.84, 16.04, 16.07, 16.04, 15.99, 15.99, 16.06, 16.16, 16.23, 16.23, 16.2, 16.15, 16.13, 16.13, 16.14, 16.15, 16.14, 16.07, 15.96, 15.82, 15.69, 15.59, 15.51, 15.44, 15.38, 15.31, 15.24, 15.14, 15.03, 14.92, 14.82, 14.73, 14.67, 14.63, 14.62, 14.61, 14.61, 14.62, 14.66, 14.71, 14.76, 14.81, 14.85, 14.89, 14.92, 14.95, 14.96, 14.96, 14.95, 14.94, 14.92, 14.89, 14.85, 14.82, 14.81, 14.81, 14.83, 14.87, 14.92, 14.95, 14.97, 14.96, 14.94, 14.9, 14.83, 14.76, 14.69, 14.63, 14.57, 14.53, 14.49, 14.46, 14.44, 14.42, 14.39, 14.38, 14.36, 14.33, 14.3, 14.25, 14.18, 14.11, 14.03, 13.96, 13.9, 13.85, 13.82, 13.83, 13.86, 13.91, 13.95, 13.98, 14.02, 14.07, 14.1, 14.13, 14.16, 14.19, 14.22, 14.26, 14.32, 14.38, 14.44, 14.52, 14.6, 14.66, 14.72, 14.77, 14.8, 14.8, 14.79, 14.77, 14.75, 14.72, 14.69, 14.66, 14.63, 14.59, 14.55, 14.5, 14.47, 14.43, 14.41, 14.38, 14.35, 14.33, 14.31, 14.29, 14.28, 14.26, 14.24, 14.23, 14.21, 14.2, 14.19, 14.18, 14.17, 14.16, 14.15, 14.13, 14.12, 14.11, 14.11, 14.1, 14.09, 14.08, 14.07, 14.06, 14.06, 14.07, 14.08, 14.1, 14.11, 14.12, 14.13, 14.14, 14.16, 14.18, 14.19, 14.22, 14.23, 14.25, 14.26, 14.27, 14.28, 14.29, 14.29, 14.3, 14.31, 14.32, 14.34, 14.35, 14.35, 14.36, 14.36, 14.34, 14.32, 14.3, 14.27, 14.25, 14.22, 14.2, 14.19, 14.18, 14.18, 14.18, 14.19, 14.19, 14.2, 14.21, 14.21, 14.22, 14.22, 14.23, 14.25, 14.27, 14.29, 14.31, 14.34, 14.36, 14.38, 14.4, 14.42, 14.44, 14.46, 14.47, 14.47, 14.48, 14.48, 14.49, 14.5, 14.5, 14.51, 14.51, 14.52, 14.52, 14.51, 14.5, 14.48, 14.46, 14.45, 14.44, 14.43, 14.43, 14.42, 14.42, 14.42, 14.42, 14.42, 14.42, 14.41, 14.41, 14.41, 14.41, 14.41, 14.42, 14.43, 14.43, 14.45, 14.45, 14.46, 14.47, 14.49, 14.5, 14.52, 14.54, 14.57, 14.6, 14.63, 14.65, 14.67, 14.7, 14.72, 14.74, 14.75, 14.76, 14.76, 14.76, 14.76, 14.77, 14.77, 14.78, 14.8, 14.81, 14.82, 14.83, 14.83, 14.84, 14.85, 14.86, 14.88, 14.9, 14.93, 14.95, 14.98, 15.0, 15.03, 15.05, 15.08, 15.1, 15.12, 15.14, 15.16, 15.18, 15.19, 15.2, 15.21, 15.22, 15.23, 15.24, 15.24, 15.26, 15.27, 15.29, 15.31, 15.33, 15.35, 15.38, 15.42, 15.46, 15.5, 15.53, 15.54, 15.55, 15.55, 15.55, 15.55, 15.56, 15.57, 15.59, 15.6, 15.62, 15.64, 15.65, 15.66, 15.68, 15.69, 15.71, 15.73, 15.75, 15.78, 15.8, 15.82, 15.84, 15.86, 15.88, 15.9, 15.91, 15.9, 15.88, 15.86, 15.84, 15.83, 15.8, 15.78, 15.76, 15.73, 15.71, 15.69, 15.66, 15.64, 15.61, 15.58, 15.54, 15.51, 15.49, 15.49, 15.5, 15.53, 15.55, 15.58, 15.6, 15.62, 15.63, 15.65, 15.66, 15.67, 15.69, 15.7, 15.71, 15.72, 15.73, 15.73, 15.74, 15.74, 15.74, 15.75, 15.75, 15.76, 15.76, 15.77, 15.77, 15.78, 15.79, 15.8, 16.46, 16.8, 17.34, 17.95, 18.46, 18.93, 19.35, 19.72, 20.09, 20.44, 20.85, 21.36, 22.13, 23.14, 24.19, 25.14, 25.91, 26.5, 26.94, 27.25, 27.45, 27.56, 27.61, 27.6, 27.56, 27.49, 27.39, 27.28, 27.16, 27.04, 26.91, 26.78, 26.65, 26.52, 26.39, 26.26, 26.12, 25.97, 25.82, 25.66, 25.51, 25.36, 25.21, 25.06, 24.92, 24.79, 24.66, 24.54, 24.43, 24.32, 24.22, 24.11, 24.0, 23.89, 23.78, 23.66, 23.54, 23.42, 23.31, 23.22, 23.13, 23.05, 22.98, 22.9, 22.83, 22.75, 22.67, 22.58, 22.49, 22.41, 22.31, 22.22, 22.13, 22.04, 21.95, 21.87, 21.78, 21.69, 21.6, 21.51, 21.44, 21.36, 21.3, 21.24, 21.2, 21.16, 21.14, 21.12, 21.12, 21.14, 21.17, 21.21, 21.27, 21.35}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {207.128, 207.122, 207.125, 207.129, 207.134, 207.143, 207.154, 207.166, 207.177, 207.199, 207.214, 207.211, 207.23, 207.242, 207.251, 207.262, 207.27, 207.268, 207.28, 207.291, 207.293, 207.302, 207.312, 207.318, 207.322, 207.325, 207.336, 207.337, 207.345, 207.35, 207.354, 207.367, 207.372, 207.379, 207.393, 207.393, 207.405, 207.407, 207.407, 207.424, 207.424, 207.422, 207.423, 207.421, 207.424, 207.418, 207.416, 207.417, 207.414, 207.417, 207.401, 207.39, 207.385, 207.375, 207.368, 207.356, 207.341, 207.336, 207.321, 207.312, 207.296, 207.284, 207.272, 207.262, 207.253, 207.238, 207.224, 207.215, 207.209, 207.196, 207.187, 207.172, 207.168, 207.159, 207.15, 207.135, 207.127, 207.117, 207.113, 207.099, 207.1, 207.083, 207.077, 207.073, 207.069, 207.065, 207.064, 207.058, 207.061, 207.065, 207.061, 207.066, 207.069, 207.069, 207.076, 207.084, 207.089, 207.104, 207.107, 207.111, 207.121, 207.128, 207.135, 207.152, 207.158, 207.17, 207.182, 207.191, 207.201, 207.212, 207.222, 207.226, 207.231, 207.237, 207.241, 207.251, 207.259, 207.266, 207.27, 207.284, 207.299, 207.311, 207.323, 207.319, 207.331, 207.335, 207.348, 207.357, 207.366, 207.377, 207.387, 207.393, 207.409, 207.413, 207.423, 207.428, 207.429, 207.432, 207.44, 207.447, 207.447, 207.439, 207.443, 207.435, 207.437, 207.433, 207.423, 207.42, 207.409, 207.4, 207.386, 207.375, 207.363, 207.345, 207.321, 207.306, 207.292, 207.279, 207.263, 207.245, 207.23, 207.212, 207.196, 207.172, 207.157, 207.142, 207.126, 207.11, 207.101, 207.093, 207.083, 207.074, 207.06, 207.049, 207.038, 207.035, 207.023, 207.016, 207.008, 207.009, 207.01, 207.013, 207.022, 207.025, 207.033, 207.043, 207.051, 207.066, 207.077, 207.087, 207.097, 207.104, 207.118, 207.121, 207.129, 207.142, 207.158, 207.164, 207.173, 207.187, 207.203, 207.21, 207.216, 207.232, 207.24, 207.246, 207.254, 207.264, 207.27, 207.277, 207.275, 207.28, 207.284, 207.285, 207.282, 207.284, 207.292, 207.304, 207.312, 207.323, 207.337, 207.349, 207.36, 207.374, 207.384, 207.401, 207.413, 207.426, 207.439, 207.457, 207.468, 207.483, 207.492, 207.499, 207.507, 207.516, 207.523, 207.528, 207.533, 207.537, 207.546, 207.547, 207.545, 207.544, 207.537, 207.522, 207.507, 207.498, 207.481, 207.457, 207.438, 207.42, 207.402, 207.379, 207.35, 207.325, 207.306, 207.279, 207.259, 207.234, 207.206, 207.192, 207.164, 207.148, 207.129, 207.112, 207.099, 207.091, 207.072, 207.06, 207.051, 207.043, 207.031, 207.029, 207.017, 207.013, 207.016, 207.016, 207.016, 207.027, 207.03, 207.029, 207.035, 207.049, 207.059, 207.063, 207.073, 207.088, 207.091, 207.104, 207.114, 207.117, 207.134, 207.142, 207.155, 207.17, 207.179, 207.202, 207.211, 207.227, 207.24, 207.246, 207.251, 207.264, 207.267, 207.281, 207.285, 207.29, 207.301, 207.309, 207.318, 207.318, 207.326, 207.342, 207.347, 207.356, 207.373, 207.379, 207.397, 207.41, 207.434, 207.448, 207.466, 207.476, 207.492, 207.514, 207.52, 207.532, 207.553, 207.563, 207.582, 207.601, 207.61, 207.624, 207.629, 207.633, 207.649, 207.657, 207.651, 207.646, 207.642, 207.634, 207.619, 207.604, 207.583, 207.581, 207.558, 207.531, 207.506, 207.483, 207.458, 207.436, 207.398, 207.372, 207.341, 207.311, 207.284, 207.268, 207.237, 207.214, 207.189, 207.165, 207.138, 207.124, 207.099, 207.079, 207.068, 207.05, 207.037, 207.025, 207.013, 207.007, 206.999, 206.994, 206.995, 206.996, 206.998, 207.01, 207.017, 207.027, 207.037, 207.046, 207.059, 207.072, 207.081, 207.096, 207.113, 207.129, 207.146, 207.154, 207.17, 207.186, 207.198, 207.204, 207.224, 207.238, 207.243, 207.248, 207.257, 207.27, 207.279, 207.283, 207.289, 207.295, 207.303, 207.31, 207.323, 207.325, 207.332, 207.336, 207.345, 207.351, 207.361, 207.36, 207.378, 207.395, 207.417, 207.431, 207.455, 207.474, 207.492, 207.515, 207.527, 207.546, 207.563, 207.576, 207.597, 207.618, 207.631, 207.648, 207.664, 207.677, 207.688, 207.696, 207.698, 207.714, 207.713, 207.71, 207.708, 207.7, 207.688, 207.667, 207.648, 207.633, 207.608, 207.582, 207.563, 207.529, 207.507, 207.482, 207.447, 207.419, 207.383, 207.353, 207.325, 207.294, 207.268, 207.24, 207.215, 207.19, 207.16, 207.131, 207.098, 207.08, 207.057, 207.04, 207.027, 207.018, 207.019, 207.014, 207.01, 206.998, 206.995, 207.0, 206.996, 207.004, 207.012, 207.021, 207.03, 207.045, 207.056, 207.074, 207.082, 207.099, 207.11, 207.133, 207.15, 207.163, 207.178, 207.194, 207.201, 207.214, 207.226, 207.231, 207.24, 207.249, 207.254, 207.261, 207.265, 207.268, 207.272, 207.27, 207.268, 207.274, 207.281, 207.278, 207.293, 207.298, 207.312, 207.32, 207.335, 207.344, 207.36, 207.374, 207.387, 207.404, 207.423, 207.447, 207.472, 207.494, 207.516, 207.538, 207.561, 207.58, 207.591, 207.618, 207.632, 207.65, 207.662, 207.678, 207.696, 207.705, 207.708, 207.711, 207.707, 207.706, 207.711, 207.698, 207.695, 207.684, 207.667, 207.647, 207.632, 207.611, 207.582, 207.55, 207.524, 207.494, 207.456, 207.423, 207.384, 207.353, 207.319, 207.293, 207.257, 207.228, 207.198, 207.167, 207.14, 207.119, 207.094, 207.07, 207.047, 207.033, 207.017, 207.003, 206.998, 206.984, 206.979, 206.969, 206.967, 206.971, 206.979, 206.981, 206.993, 206.999, 207.013, 207.022, 207.037, 207.056, 207.065, 207.092, 207.106, 207.117, 207.145, 207.159, 207.179, 207.201, 207.215, 207.23, 207.239, 195.962, 0.585, 0.586, 0.579, 0.571, 0.569, 0.561, 0.557, 0.549, 0.539, 0.536, 0.524, 0.497, 0.488, 0.477, 0.465, 0.451, 0.439, 0.425, 0.42, 0.412, 0.41, 0.406, 0.402, 0.403, 0.401, 0.402, 0.404, 0.405, 0.41, 0.409, 0.413, 0.414, 0.421, 0.42, 0.423, 0.428, 0.433, 0.434, 0.439, 0.442, 0.441, 0.443, 0.445, 0.451, 0.45, 0.456, 0.457, 0.458, 0.457, 0.46, 0.463, 0.464, 0.468, 0.47, 0.474, 0.474, 0.477, 0.476, 0.478, 0.481, 0.478, 0.479, 0.483, 0.483, 0.484, 0.485, 0.487, 0.485, 0.489, 0.492, 0.495, 0.496, 0.501, 0.502, 0.506, 0.505, 0.508, 0.506, 0.511, 0.51, 0.515, 0.515, 0.518, 0.519, 0.525, 0.525, 0.526, 0.526, 0.524, 0.528, 0.523, 0.526, 0.524, 0.526}
PRES_REL_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {205.58421, 205.58456, 205.58444, 205.58757, 205.59082, 205.59721, 205.61368, 205.62344, 205.64, 205.65588, 205.67235, 205.67252, 205.69215, 205.69835, 205.70474, 205.72127, 205.72438, 205.721, 205.73755, 205.74725, 205.7471, 205.76384, 205.76672, 205.77325, 205.77997, 205.77979, 205.79625, 205.79282, 205.8027, 205.80595, 205.8091, 205.82217, 205.83221, 205.8352, 205.84473, 205.84473, 205.86142, 205.86461, 205.86461, 205.88097, 205.88097, 205.87761, 205.88097, 205.88112, 205.88097, 205.87091, 205.871, 205.87442, 205.86775, 205.87442, 205.8547, 205.8449, 205.84523, 205.83203, 205.82555, 205.81241, 205.79959, 205.79625, 205.7731, 205.76672, 205.75383, 205.74074, 205.72763, 205.72127, 205.70808, 205.69513, 205.68561, 205.66884, 205.66911, 205.64922, 205.64291, 205.62999, 205.62329, 205.61691, 205.61052, 205.59406, 205.58766, 205.5745, 205.57129, 205.55821, 205.55821, 205.54202, 205.53548, 205.52885, 205.53238, 205.52568, 205.5224, 205.51587, 205.52255, 205.52568, 205.52255, 205.52568, 205.53238, 205.53238, 205.53548, 205.54532, 205.54857, 205.56143, 205.56131, 205.56798, 205.57768, 205.58421, 205.59406, 205.61389, 205.62038, 205.62665, 205.63966, 205.64955, 205.65932, 205.66902, 205.6822, 205.6854, 205.68864, 205.69513, 205.70183, 205.70474, 205.71463, 205.72797, 205.72438, 205.74074, 205.75711, 205.77017, 205.77641, 205.78006, 205.78633, 205.79298, 205.80255, 205.8089, 205.82567, 205.83542, 205.84506, 205.84473, 205.86452, 205.87122, 205.88097, 205.88416, 205.88069, 205.89078, 205.89723, 205.90372, 205.90372, 205.89386, 205.89703, 205.89064, 205.89055, 205.88731, 205.88097, 205.87424, 205.86452, 205.85812, 205.8418, 205.83203, 205.81895, 205.8027, 205.7731, 205.76018, 205.75058, 205.73755, 205.72127, 205.70502, 205.69215, 205.66902, 205.64922, 205.62999, 205.61356, 205.60066, 205.5809, 205.56798, 205.56158, 205.55167, 205.54202, 205.5321, 205.51576, 205.50597, 205.49623, 205.49644, 205.48335, 205.4803, 205.47046, 205.46696, 205.47023, 205.47012, 205.47998, 205.48668, 205.49657, 205.49942, 205.50938, 205.52568, 205.53548, 205.54518, 205.55846, 205.56143, 205.57784, 205.57768, 205.58757, 205.60066, 205.62038, 205.62004, 205.6333, 205.64291, 205.66257, 205.66565, 205.67566, 205.68518, 205.695, 205.70149, 205.71138, 205.72466, 205.72438, 205.73772, 205.73434, 205.73755, 205.74074, 205.7407, 205.7374, 205.74074, 205.75058, 205.75684, 205.76672, 205.77641, 205.79282, 205.80939, 205.81914, 205.82867, 205.83836, 205.8547, 205.87122, 205.88077, 205.89386, 205.91696, 205.92668, 205.93959, 205.94598, 205.95245, 205.96234, 205.97559, 205.97859, 205.98184, 205.9918, 205.98824, 206.00494, 206.00148, 205.99806, 206.0016, 205.98824, 205.97531, 205.96234, 205.95245, 205.93625, 205.91696, 205.89732, 205.87424, 205.86151, 205.8352, 205.80595, 205.77979, 205.76018, 205.73755, 205.71463, 205.68848, 205.66249, 205.65292, 205.62004, 205.60713, 205.58757, 205.57129, 205.55821, 205.55185, 205.53229, 205.51576, 205.50938, 205.49942, 205.49323, 205.48984, 205.47682, 205.47012, 205.4803, 205.4803, 205.4803, 205.48653, 205.48984, 205.48984, 205.49644, 205.50597, 205.5192, 205.5224, 205.52885, 205.54857, 205.55185, 205.56143, 205.57463, 205.5745, 205.59082, 205.60066, 205.61368, 205.62665, 205.63303, 205.65929, 205.67252, 205.68536, 205.695, 205.70149, 205.70474, 205.72466, 205.72453, 205.74083, 205.7407, 205.74728, 205.75696, 205.76685, 205.77325, 205.77325, 205.78308, 205.79604, 205.80608, 205.81241, 205.82872, 205.8352, 205.85144, 205.86452, 205.89064, 205.90024, 205.92331, 205.93304, 205.94598, 205.97226, 205.97198, 205.98851, 206.00789, 206.02116, 206.04076, 206.05695, 206.06677, 206.0763, 206.0864, 206.08957, 206.1024, 206.11238, 206.10225, 206.10258, 206.0959, 206.08606, 206.07312, 206.0602, 206.03732, 206.03387, 206.01115, 205.98851, 205.96234, 205.93959, 205.91348, 205.89404, 205.85481, 205.83221, 205.79959, 205.77017, 205.74074, 205.721, 205.69513, 205.67235, 205.64627, 205.62344, 205.59746, 205.57759, 205.55821, 205.53539, 205.52556, 205.51285, 205.49295, 205.48668, 205.47012, 205.46358, 205.46051, 205.45404, 205.45741, 205.45393, 205.45723, 205.47023, 205.47682, 205.48653, 205.49295, 205.50615, 205.5192, 205.53229, 205.53865, 205.55157, 205.57129, 205.58757, 205.60385, 205.61368, 205.62665, 205.64638, 205.65265, 205.6591, 205.68561, 205.69513, 205.70168, 205.7049, 205.71129, 205.72438, 205.73755, 205.74426, 205.74393, 205.75047, 205.76036, 205.76682, 205.77641, 205.77979, 205.78961, 205.79625, 205.8027, 205.80917, 205.8156, 205.81914, 205.83188, 205.84816, 205.87442, 205.884, 205.91367, 205.93317, 205.94598, 205.96877, 205.98532, 206.00494, 206.02116, 206.03078, 206.05368, 206.07663, 206.08615, 206.10243, 206.11534, 206.1284, 206.145, 206.14798, 206.14789, 206.1676, 206.16429, 206.16447, 206.16106, 206.1512, 206.145, 206.122, 206.10243, 206.08957, 206.06343, 206.04076, 206.02116, 205.98514, 205.96234, 205.93625, 205.90372, 205.8777, 205.84189, 205.81259, 205.77979, 205.75398, 205.721, 205.695, 205.66884, 205.64955, 205.6134, 205.59093, 205.55496, 205.54218, 205.51587, 205.49962, 205.48653, 205.47333, 205.48013, 205.47694, 205.47023, 205.45723, 205.45741, 205.46051, 205.45393, 205.46375, 205.4736, 205.47998, 205.48984, 205.50284, 205.51251, 205.5321, 205.54202, 205.55821, 205.56798, 205.59427, 205.61052, 205.62354, 205.63652, 205.65622, 205.65932, 205.67235, 205.6854, 205.68864, 205.695, 205.7049, 205.71138, 205.71799, 205.72108, 205.721, 205.72763, 205.72438, 205.721, 205.731, 205.74083, 205.73418, 205.7471, 205.75711, 205.76672, 205.77654, 205.79298, 205.79936, 205.81914, 205.82867, 205.84506, 205.86142, 205.88097, 205.90372, 205.92986, 205.94933, 205.97559, 205.99512, 206.01779, 206.0374, 206.04713, 206.07663, 206.08615, 206.10577, 206.11205, 206.13176, 206.14798, 206.16125, 206.16106, 206.16779, 206.16457, 206.15778, 206.16779, 206.14789, 206.14798, 206.13837, 206.122, 206.09915, 206.08615, 206.06331, 206.04076, 206.00809, 205.97859, 205.94933, 205.91016, 205.88097, 205.83836, 205.81259, 205.78006, 205.7471, 205.71129, 205.68875, 205.65265, 205.62677, 205.5973, 205.57784, 205.55167, 205.52893, 205.50615, 205.49657, 205.47682, 205.46033, 205.45723, 205.44077, 205.43759, 205.42793, 205.42453, 205.42773, 205.43759, 205.44101, 205.45404, 205.46051, 205.47012, 205.47998, 205.49295, 205.51251, 205.52568, 205.54842, 205.56482, 205.5745, 205.60048, 205.61691, 205.63303, 205.65932, 205.66884, 205.69215, 205.69855, 194.51114, 0.58396745, 0.58050436, 0.5736349, 0.5633157, 0.56332886, 0.5599226, 0.5530342, 0.54271483, 0.5324089, 0.5324278, 0.52213305, 0.49465123, 0.48433733, 0.47403675, 0.46028638, 0.4500046, 0.43625405, 0.42251462, 0.41563377, 0.41222718, 0.40878293, 0.40535197, 0.39846346, 0.40191314, 0.40192652, 0.39846346, 0.40190756, 0.3984445, 0.40878293, 0.40533298, 0.4087641, 0.412214, 0.41908374, 0.41563377, 0.42252797, 0.42595348, 0.42592144, 0.43282866, 0.43625405, 0.44314831, 0.43624085, 0.43968517, 0.44312933, 0.4500046, 0.4465547, 0.45343003, 0.45687985, 0.45341685, 0.45687985, 0.45686096, 0.45684218, 0.4637495, 0.46718055, 0.47062477, 0.46714288, 0.46714288, 0.47403675, 0.4705871, 0.47403118, 0.48092535, 0.47403118, 0.47748098, 0.48436955, 0.48436955, 0.4809064, 0.47744346, 0.4808875, 0.47744346, 0.48433173, 0.49122575, 0.49120697, 0.49465677, 0.49808225, 0.4946191, 0.5015076, 0.50497055, 0.5049518, 0.5015076, 0.51184595, 0.5049385, 0.5083638, 0.5083638, 0.5152579, 0.51525235, 0.52212745, 0.52212745, 0.51866436, 0.51866436, 0.52213305, 0.5221083, 0.51868325, 0.51866436, 0.52213305, 0.51866436}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
