netcdf file-160.nc {
  dimensions:
    DEPTH = 25;
  variables:
    float LATITUDE(DEPTH=25);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=25);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=25);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=25);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=25);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=25);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222, 22383.065659722222}
TEMP =
  {26.4149, 26.3853, 26.3546, 26.3282, 26.3097, 26.2955, 26.2955, 26.2994, 26.3077, 26.3217, 26.3324, 26.3343, 26.3306, 26.3244, 26.3192, 26.3252, 26.3646, 26.4219, 26.441, 26.4486, 26.4579, 26.4742, 26.4997, 26.5155, 26.5272}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.908, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841}
}
