netcdf IMOS_ANMN-TS_20150113T230000Z_WATR20_FV01_WATR20-1407-Seabird-SBE39-600m-temp-press.-25_END-20150122T025000Z_id-7734.nc {
  dimensions:
    TIME = UNLIMITED;   // (1176 currently)
  variables:
    double TIME(TIME=1176);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=1176);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=1176);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=1176);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=1176);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=1176);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=1176);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=1176);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=1176);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=1176);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=1176);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=1176);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=1176);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :instrument = "Seabird         SBE39 [600m] temp & press.";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "3949303-4207";
  :history = "2015-01-29T06:32:02Z - depthPP: Depth computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and relative pressure measurements (calibration offset usually performed to balance current atmospheric pressure and acute sensor precision at a deployed depth).";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 25.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = -0.285143f; // float
  :geospatial_vertical_max = 35.716064f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-22T02:50:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.965277777777, 23753.972222222223, 23753.979166666668, 23753.98611111111, 23753.993055555555, 23754.0, 23754.006944444445, 23754.01388888889, 23754.020833333332, 23754.027777777777, 23754.034722222223, 23754.041666666668, 23754.04861111111, 23754.055555555555, 23754.0625, 23754.069444444445, 23754.07638888889, 23754.083333333332, 23754.090277777777, 23754.097222222223, 23754.104166666668, 23754.11111111111, 23754.118055555555, 23754.125, 23754.131944444445, 23754.13888888889, 23754.145833333332, 23754.152777777777, 23754.159722222223, 23754.166666666668, 23754.17361111111, 23754.180555555555, 23754.1875, 23754.194444444445, 23754.20138888889, 23754.208333333332, 23754.215277777777, 23754.222222222223, 23754.229166666668, 23754.23611111111, 23754.243055555555, 23754.25, 23754.256944444445, 23754.26388888889, 23754.270833333332, 23754.277777777777, 23754.284722222223, 23754.291666666668, 23754.29861111111, 23754.305555555555, 23754.3125, 23754.319444444445, 23754.32638888889, 23754.333333333332, 23754.340277777777, 23754.347222222223, 23754.354166666668, 23754.36111111111, 23754.368055555555, 23754.375, 23754.381944444445, 23754.38888888889, 23754.395833333332, 23754.402777777777, 23754.409722222223, 23754.416666666668, 23754.42361111111, 23754.430555555555, 23754.4375, 23754.444444444445, 23754.45138888889, 23754.458333333332, 23754.465277777777, 23754.472222222223, 23754.479166666668, 23754.48611111111, 23754.493055555555, 23754.5, 23754.506944444445, 23754.51388888889, 23754.520833333332, 23754.527777777777, 23754.534722222223, 23754.541666666668, 23754.54861111111, 23754.555555555555, 23754.5625, 23754.569444444445, 23754.57638888889, 23754.583333333332, 23754.590277777777, 23754.597222222223, 23754.604166666668, 23754.61111111111, 23754.618055555555, 23754.625, 23754.631944444445, 23754.63888888889, 23754.645833333332, 23754.652777777777, 23754.659722222223, 23754.666666666668, 23754.67361111111, 23754.680555555555, 23754.6875, 23754.694444444445, 23754.70138888889, 23754.708333333332, 23754.715277777777, 23754.722222222223, 23754.729166666668, 23754.73611111111, 23754.743055555555, 23754.75, 23754.756944444445, 23754.76388888889, 23754.770833333332, 23754.777777777777, 23754.784722222223, 23754.791666666668, 23754.79861111111, 23754.805555555555, 23754.8125, 23754.819444444445, 23754.82638888889, 23754.833333333332, 23754.840277777777, 23754.847222222223, 23754.854166666668, 23754.86111111111, 23754.868055555555, 23754.875, 23754.881944444445, 23754.88888888889, 23754.895833333332, 23754.902777777777, 23754.909722222223, 23754.916666666668, 23754.92361111111, 23754.930555555555, 23754.9375, 23754.944444444445, 23754.95138888889, 23754.958333333332, 23754.965277777777, 23754.972222222223, 23754.979166666668, 23754.98611111111, 23754.993055555555, 23755.0, 23755.006944444445, 23755.01388888889, 23755.020833333332, 23755.027777777777, 23755.034722222223, 23755.041666666668, 23755.04861111111, 23755.055555555555, 23755.0625, 23755.069444444445, 23755.07638888889, 23755.083333333332, 23755.090277777777, 23755.097222222223, 23755.104166666668, 23755.11111111111, 23755.118055555555, 23755.125, 23755.131944444445, 23755.13888888889, 23755.145833333332, 23755.152777777777, 23755.159722222223, 23755.166666666668, 23755.17361111111, 23755.180555555555, 23755.1875, 23755.194444444445, 23755.20138888889, 23755.208333333332, 23755.215277777777, 23755.222222222223, 23755.229166666668, 23755.23611111111, 23755.243055555555, 23755.25, 23755.256944444445, 23755.26388888889, 23755.270833333332, 23755.277777777777, 23755.284722222223, 23755.291666666668, 23755.29861111111, 23755.305555555555, 23755.3125, 23755.319444444445, 23755.32638888889, 23755.333333333332, 23755.340277777777, 23755.347222222223, 23755.354166666668, 23755.36111111111, 23755.368055555555, 23755.375, 23755.381944444445, 23755.38888888889, 23755.395833333332, 23755.402777777777, 23755.409722222223, 23755.416666666668, 23755.42361111111, 23755.430555555555, 23755.4375, 23755.444444444445, 23755.45138888889, 23755.458333333332, 23755.465277777777, 23755.472222222223, 23755.479166666668, 23755.48611111111, 23755.493055555555, 23755.5, 23755.506944444445, 23755.51388888889, 23755.520833333332, 23755.527777777777, 23755.534722222223, 23755.541666666668, 23755.54861111111, 23755.555555555555, 23755.5625, 23755.569444444445, 23755.57638888889, 23755.583333333332, 23755.590277777777, 23755.597222222223, 23755.604166666668, 23755.61111111111, 23755.618055555555, 23755.625, 23755.631944444445, 23755.63888888889, 23755.645833333332, 23755.652777777777, 23755.659722222223, 23755.666666666668, 23755.67361111111, 23755.680555555555, 23755.6875, 23755.694444444445, 23755.70138888889, 23755.708333333332, 23755.715277777777, 23755.722222222223, 23755.729166666668, 23755.73611111111, 23755.743055555555, 23755.75, 23755.756944444445, 23755.76388888889, 23755.770833333332, 23755.777777777777, 23755.784722222223, 23755.791666666668, 23755.79861111111, 23755.805555555555, 23755.8125, 23755.819444444445, 23755.82638888889, 23755.833333333332, 23755.840277777777, 23755.847222222223, 23755.854166666668, 23755.86111111111, 23755.868055555555, 23755.875, 23755.881944444445, 23755.88888888889, 23755.895833333332, 23755.902777777777, 23755.909722222223, 23755.916666666668, 23755.92361111111, 23755.930555555555, 23755.9375, 23755.944444444445, 23755.95138888889, 23755.958333333332, 23755.965277777777, 23755.972222222223, 23755.979166666668, 23755.98611111111, 23755.993055555555, 23756.0, 23756.006944444445, 23756.01388888889, 23756.020833333332, 23756.027777777777, 23756.034722222223, 23756.041666666668, 23756.04861111111, 23756.055555555555, 23756.0625, 23756.069444444445, 23756.07638888889, 23756.083333333332, 23756.090277777777, 23756.097222222223, 23756.104166666668, 23756.11111111111, 23756.118055555555, 23756.125, 23756.131944444445, 23756.13888888889, 23756.145833333332, 23756.152777777777, 23756.159722222223, 23756.166666666668, 23756.17361111111, 23756.180555555555, 23756.1875, 23756.194444444445, 23756.20138888889, 23756.208333333332, 23756.215277777777, 23756.222222222223, 23756.229166666668, 23756.23611111111, 23756.243055555555, 23756.25, 23756.256944444445, 23756.26388888889, 23756.270833333332, 23756.277777777777, 23756.284722222223, 23756.291666666668, 23756.29861111111, 23756.305555555555, 23756.3125, 23756.319444444445, 23756.32638888889, 23756.333333333332, 23756.340277777777, 23756.347222222223, 23756.354166666668, 23756.36111111111, 23756.368055555555, 23756.375, 23756.381944444445, 23756.38888888889, 23756.395833333332, 23756.402777777777, 23756.409722222223, 23756.416666666668, 23756.42361111111, 23756.430555555555, 23756.4375, 23756.444444444445, 23756.45138888889, 23756.458333333332, 23756.465277777777, 23756.472222222223, 23756.479166666668, 23756.48611111111, 23756.493055555555, 23756.5, 23756.506944444445, 23756.51388888889, 23756.520833333332, 23756.527777777777, 23756.534722222223, 23756.541666666668, 23756.54861111111, 23756.555555555555, 23756.5625, 23756.569444444445, 23756.57638888889, 23756.583333333332, 23756.590277777777, 23756.597222222223, 23756.604166666668, 23756.61111111111, 23756.618055555555, 23756.625, 23756.631944444445, 23756.63888888889, 23756.645833333332, 23756.652777777777, 23756.659722222223, 23756.666666666668, 23756.67361111111, 23756.680555555555, 23756.6875, 23756.694444444445, 23756.70138888889, 23756.708333333332, 23756.715277777777, 23756.722222222223, 23756.729166666668, 23756.73611111111, 23756.743055555555, 23756.75, 23756.756944444445, 23756.76388888889, 23756.770833333332, 23756.777777777777, 23756.784722222223, 23756.791666666668, 23756.79861111111, 23756.805555555555, 23756.8125, 23756.819444444445, 23756.82638888889, 23756.833333333332, 23756.840277777777, 23756.847222222223, 23756.854166666668, 23756.86111111111, 23756.868055555555, 23756.875, 23756.881944444445, 23756.88888888889, 23756.895833333332, 23756.902777777777, 23756.909722222223, 23756.916666666668, 23756.92361111111, 23756.930555555555, 23756.9375, 23756.944444444445, 23756.95138888889, 23756.958333333332, 23756.965277777777, 23756.972222222223, 23756.979166666668, 23756.98611111111, 23756.993055555555, 23757.0, 23757.006944444445, 23757.01388888889, 23757.020833333332, 23757.027777777777, 23757.034722222223, 23757.041666666668, 23757.04861111111, 23757.055555555555, 23757.0625, 23757.069444444445, 23757.07638888889, 23757.083333333332, 23757.090277777777, 23757.097222222223, 23757.104166666668, 23757.11111111111, 23757.118055555555, 23757.125, 23757.131944444445, 23757.13888888889, 23757.145833333332, 23757.152777777777, 23757.159722222223, 23757.166666666668, 23757.17361111111, 23757.180555555555, 23757.1875, 23757.194444444445, 23757.20138888889, 23757.208333333332, 23757.215277777777, 23757.222222222223, 23757.229166666668, 23757.23611111111, 23757.243055555555, 23757.25, 23757.256944444445, 23757.26388888889, 23757.270833333332, 23757.277777777777, 23757.284722222223, 23757.291666666668, 23757.29861111111, 23757.305555555555, 23757.3125, 23757.319444444445, 23757.32638888889, 23757.333333333332, 23757.340277777777, 23757.347222222223, 23757.354166666668, 23757.36111111111, 23757.368055555555, 23757.375, 23757.381944444445, 23757.38888888889, 23757.395833333332, 23757.402777777777, 23757.409722222223, 23757.416666666668, 23757.42361111111, 23757.430555555555, 23757.4375, 23757.444444444445, 23757.45138888889, 23757.458333333332, 23757.465277777777, 23757.472222222223, 23757.479166666668, 23757.48611111111, 23757.493055555555, 23757.5, 23757.506944444445, 23757.51388888889, 23757.520833333332, 23757.527777777777, 23757.534722222223, 23757.541666666668, 23757.54861111111, 23757.555555555555, 23757.5625, 23757.569444444445, 23757.57638888889, 23757.583333333332, 23757.590277777777, 23757.597222222223, 23757.604166666668, 23757.61111111111, 23757.618055555555, 23757.625, 23757.631944444445, 23757.63888888889, 23757.645833333332, 23757.652777777777, 23757.659722222223, 23757.666666666668, 23757.67361111111, 23757.680555555555, 23757.6875, 23757.694444444445, 23757.70138888889, 23757.708333333332, 23757.715277777777, 23757.722222222223, 23757.729166666668, 23757.73611111111, 23757.743055555555, 23757.75, 23757.756944444445, 23757.76388888889, 23757.770833333332, 23757.777777777777, 23757.784722222223, 23757.791666666668, 23757.79861111111, 23757.805555555555, 23757.8125, 23757.819444444445, 23757.82638888889, 23757.833333333332, 23757.840277777777, 23757.847222222223, 23757.854166666668, 23757.86111111111, 23757.868055555555, 23757.875, 23757.881944444445, 23757.88888888889, 23757.895833333332, 23757.902777777777, 23757.909722222223, 23757.916666666668, 23757.92361111111, 23757.930555555555, 23757.9375, 23757.944444444445, 23757.95138888889, 23757.958333333332, 23757.965277777777, 23757.972222222223, 23757.979166666668, 23757.98611111111, 23757.993055555555, 23758.0, 23758.006944444445, 23758.01388888889, 23758.020833333332, 23758.027777777777, 23758.034722222223, 23758.041666666668, 23758.04861111111, 23758.055555555555, 23758.0625, 23758.069444444445, 23758.07638888889, 23758.083333333332, 23758.090277777777, 23758.097222222223, 23758.104166666668, 23758.11111111111, 23758.118055555555, 23758.125, 23758.131944444445, 23758.13888888889, 23758.145833333332, 23758.152777777777, 23758.159722222223, 23758.166666666668, 23758.17361111111, 23758.180555555555, 23758.1875, 23758.194444444445, 23758.20138888889, 23758.208333333332, 23758.215277777777, 23758.222222222223, 23758.229166666668, 23758.23611111111, 23758.243055555555, 23758.25, 23758.256944444445, 23758.26388888889, 23758.270833333332, 23758.277777777777, 23758.284722222223, 23758.291666666668, 23758.29861111111, 23758.305555555555, 23758.3125, 23758.319444444445, 23758.32638888889, 23758.333333333332, 23758.340277777777, 23758.347222222223, 23758.354166666668, 23758.36111111111, 23758.368055555555, 23758.375, 23758.381944444445, 23758.38888888889, 23758.395833333332, 23758.402777777777, 23758.409722222223, 23758.416666666668, 23758.42361111111, 23758.430555555555, 23758.4375, 23758.444444444445, 23758.45138888889, 23758.458333333332, 23758.465277777777, 23758.472222222223, 23758.479166666668, 23758.48611111111, 23758.493055555555, 23758.5, 23758.506944444445, 23758.51388888889, 23758.520833333332, 23758.527777777777, 23758.534722222223, 23758.541666666668, 23758.54861111111, 23758.555555555555, 23758.5625, 23758.569444444445, 23758.57638888889, 23758.583333333332, 23758.590277777777, 23758.597222222223, 23758.604166666668, 23758.61111111111, 23758.618055555555, 23758.625, 23758.631944444445, 23758.63888888889, 23758.645833333332, 23758.652777777777, 23758.659722222223, 23758.666666666668, 23758.67361111111, 23758.680555555555, 23758.6875, 23758.694444444445, 23758.70138888889, 23758.708333333332, 23758.715277777777, 23758.722222222223, 23758.729166666668, 23758.73611111111, 23758.743055555555, 23758.75, 23758.756944444445, 23758.76388888889, 23758.770833333332, 23758.777777777777, 23758.784722222223, 23758.791666666668, 23758.79861111111, 23758.805555555555, 23758.8125, 23758.819444444445, 23758.82638888889, 23758.833333333332, 23758.840277777777, 23758.847222222223, 23758.854166666668, 23758.86111111111, 23758.868055555555, 23758.875, 23758.881944444445, 23758.88888888889, 23758.895833333332, 23758.902777777777, 23758.909722222223, 23758.916666666668, 23758.92361111111, 23758.930555555555, 23758.9375, 23758.944444444445, 23758.95138888889, 23758.958333333332, 23758.965277777777, 23758.972222222223, 23758.979166666668, 23758.98611111111, 23758.993055555555, 23759.0, 23759.006944444445, 23759.01388888889, 23759.020833333332, 23759.027777777777, 23759.034722222223, 23759.041666666668, 23759.04861111111, 23759.055555555555, 23759.0625, 23759.069444444445, 23759.07638888889, 23759.083333333332, 23759.090277777777, 23759.097222222223, 23759.104166666668, 23759.11111111111, 23759.118055555555, 23759.125, 23759.131944444445, 23759.13888888889, 23759.145833333332, 23759.152777777777, 23759.159722222223, 23759.166666666668, 23759.17361111111, 23759.180555555555, 23759.1875, 23759.194444444445, 23759.20138888889, 23759.208333333332, 23759.215277777777, 23759.222222222223, 23759.229166666668, 23759.23611111111, 23759.243055555555, 23759.25, 23759.256944444445, 23759.26388888889, 23759.270833333332, 23759.277777777777, 23759.284722222223, 23759.291666666668, 23759.29861111111, 23759.305555555555, 23759.3125, 23759.319444444445, 23759.32638888889, 23759.333333333332, 23759.340277777777, 23759.347222222223, 23759.354166666668, 23759.36111111111, 23759.368055555555, 23759.375, 23759.381944444445, 23759.38888888889, 23759.395833333332, 23759.402777777777, 23759.409722222223, 23759.416666666668, 23759.42361111111, 23759.430555555555, 23759.4375, 23759.444444444445, 23759.45138888889, 23759.458333333332, 23759.465277777777, 23759.472222222223, 23759.479166666668, 23759.48611111111, 23759.493055555555, 23759.5, 23759.506944444445, 23759.51388888889, 23759.520833333332, 23759.527777777777, 23759.534722222223, 23759.541666666668, 23759.54861111111, 23759.555555555555, 23759.5625, 23759.569444444445, 23759.57638888889, 23759.583333333332, 23759.590277777777, 23759.597222222223, 23759.604166666668, 23759.61111111111, 23759.618055555555, 23759.625, 23759.631944444445, 23759.63888888889, 23759.645833333332, 23759.652777777777, 23759.659722222223, 23759.666666666668, 23759.67361111111, 23759.680555555555, 23759.6875, 23759.694444444445, 23759.70138888889, 23759.708333333332, 23759.715277777777, 23759.722222222223, 23759.729166666668, 23759.73611111111, 23759.743055555555, 23759.75, 23759.756944444445, 23759.76388888889, 23759.770833333332, 23759.777777777777, 23759.784722222223, 23759.791666666668, 23759.79861111111, 23759.805555555555, 23759.8125, 23759.819444444445, 23759.82638888889, 23759.833333333332, 23759.840277777777, 23759.847222222223, 23759.854166666668, 23759.86111111111, 23759.868055555555, 23759.875, 23759.881944444445, 23759.88888888889, 23759.895833333332, 23759.902777777777, 23759.909722222223, 23759.916666666668, 23759.92361111111, 23759.930555555555, 23759.9375, 23759.944444444445, 23759.95138888889, 23759.958333333332, 23759.965277777777, 23759.972222222223, 23759.979166666668, 23759.98611111111, 23759.993055555555, 23760.0, 23760.006944444445, 23760.01388888889, 23760.020833333332, 23760.027777777777, 23760.034722222223, 23760.041666666668, 23760.04861111111, 23760.055555555555, 23760.0625, 23760.069444444445, 23760.07638888889, 23760.083333333332, 23760.090277777777, 23760.097222222223, 23760.104166666668, 23760.11111111111, 23760.118055555555, 23760.125, 23760.131944444445, 23760.13888888889, 23760.145833333332, 23760.152777777777, 23760.159722222223, 23760.166666666668, 23760.17361111111, 23760.180555555555, 23760.1875, 23760.194444444445, 23760.20138888889, 23760.208333333332, 23760.215277777777, 23760.222222222223, 23760.229166666668, 23760.23611111111, 23760.243055555555, 23760.25, 23760.256944444445, 23760.26388888889, 23760.270833333332, 23760.277777777777, 23760.284722222223, 23760.291666666668, 23760.29861111111, 23760.305555555555, 23760.3125, 23760.319444444445, 23760.32638888889, 23760.333333333332, 23760.340277777777, 23760.347222222223, 23760.354166666668, 23760.36111111111, 23760.368055555555, 23760.375, 23760.381944444445, 23760.38888888889, 23760.395833333332, 23760.402777777777, 23760.409722222223, 23760.416666666668, 23760.42361111111, 23760.430555555555, 23760.4375, 23760.444444444445, 23760.45138888889, 23760.458333333332, 23760.465277777777, 23760.472222222223, 23760.479166666668, 23760.48611111111, 23760.493055555555, 23760.5, 23760.506944444445, 23760.51388888889, 23760.520833333332, 23760.527777777777, 23760.534722222223, 23760.541666666668, 23760.54861111111, 23760.555555555555, 23760.5625, 23760.569444444445, 23760.57638888889, 23760.583333333332, 23760.590277777777, 23760.597222222223, 23760.604166666668, 23760.61111111111, 23760.618055555555, 23760.625, 23760.631944444445, 23760.63888888889, 23760.645833333332, 23760.652777777777, 23760.659722222223, 23760.666666666668, 23760.67361111111, 23760.680555555555, 23760.6875, 23760.694444444445, 23760.70138888889, 23760.708333333332, 23760.715277777777, 23760.722222222223, 23760.729166666668, 23760.73611111111, 23760.743055555555, 23760.75, 23760.756944444445, 23760.76388888889, 23760.770833333332, 23760.777777777777, 23760.784722222223, 23760.791666666668, 23760.79861111111, 23760.805555555555, 23760.8125, 23760.819444444445, 23760.82638888889, 23760.833333333332, 23760.840277777777, 23760.847222222223, 23760.854166666668, 23760.86111111111, 23760.868055555555, 23760.875, 23760.881944444445, 23760.88888888889, 23760.895833333332, 23760.902777777777, 23760.909722222223, 23760.916666666668, 23760.92361111111, 23760.930555555555, 23760.9375, 23760.944444444445, 23760.95138888889, 23760.958333333332, 23760.965277777777, 23760.972222222223, 23760.979166666668, 23760.98611111111, 23760.993055555555, 23761.0, 23761.006944444445, 23761.01388888889, 23761.020833333332, 23761.027777777777, 23761.034722222223, 23761.041666666668, 23761.04861111111, 23761.055555555555, 23761.0625, 23761.069444444445, 23761.07638888889, 23761.083333333332, 23761.090277777777, 23761.097222222223, 23761.104166666668, 23761.11111111111, 23761.118055555555, 23761.125, 23761.131944444445, 23761.13888888889, 23761.145833333332, 23761.152777777777, 23761.159722222223, 23761.166666666668, 23761.17361111111, 23761.180555555555, 23761.1875, 23761.194444444445, 23761.20138888889, 23761.208333333332, 23761.215277777777, 23761.222222222223, 23761.229166666668, 23761.23611111111, 23761.243055555555, 23761.25, 23761.256944444445, 23761.26388888889, 23761.270833333332, 23761.277777777777, 23761.284722222223, 23761.291666666668, 23761.29861111111, 23761.305555555555, 23761.3125, 23761.319444444445, 23761.32638888889, 23761.333333333332, 23761.340277777777, 23761.347222222223, 23761.354166666668, 23761.36111111111, 23761.368055555555, 23761.375, 23761.381944444445, 23761.38888888889, 23761.395833333332, 23761.402777777777, 23761.409722222223, 23761.416666666668, 23761.42361111111, 23761.430555555555, 23761.4375, 23761.444444444445, 23761.45138888889, 23761.458333333332, 23761.465277777777, 23761.472222222223, 23761.479166666668, 23761.48611111111, 23761.493055555555, 23761.5, 23761.506944444445, 23761.51388888889, 23761.520833333332, 23761.527777777777, 23761.534722222223, 23761.541666666668, 23761.54861111111, 23761.555555555555, 23761.5625, 23761.569444444445, 23761.57638888889, 23761.583333333332, 23761.590277777777, 23761.597222222223, 23761.604166666668, 23761.61111111111, 23761.618055555555, 23761.625, 23761.631944444445, 23761.63888888889, 23761.645833333332, 23761.652777777777, 23761.659722222223, 23761.666666666668, 23761.67361111111, 23761.680555555555, 23761.6875, 23761.694444444445, 23761.70138888889, 23761.708333333332, 23761.715277777777, 23761.722222222223, 23761.729166666668, 23761.73611111111, 23761.743055555555, 23761.75, 23761.756944444445, 23761.76388888889, 23761.770833333332, 23761.777777777777, 23761.784722222223, 23761.791666666668, 23761.79861111111, 23761.805555555555, 23761.8125, 23761.819444444445, 23761.82638888889, 23761.833333333332, 23761.840277777777, 23761.847222222223, 23761.854166666668, 23761.86111111111, 23761.868055555555, 23761.875, 23761.881944444445, 23761.88888888889, 23761.895833333332, 23761.902777777777, 23761.909722222223, 23761.916666666668, 23761.92361111111, 23761.930555555555, 23761.9375, 23761.944444444445, 23761.95138888889, 23761.958333333332, 23761.965277777777, 23761.972222222223, 23761.979166666668, 23761.98611111111, 23761.993055555555, 23762.0, 23762.006944444445, 23762.01388888889, 23762.020833333332, 23762.027777777777, 23762.034722222223, 23762.041666666668, 23762.04861111111, 23762.055555555555, 23762.0625, 23762.069444444445, 23762.07638888889, 23762.083333333332, 23762.090277777777, 23762.097222222223, 23762.104166666668, 23762.11111111111, 23762.118055555555}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =25.0
TEMP =
  {20.6362, 20.6409, 20.6319, 20.6585, 20.675, 20.6792, 20.742, 20.8593, 20.5804, 20.6322, 20.6389, 20.621, 20.6057, 20.5564, 20.5859, 20.7829, 20.7022, 20.6894, 20.6143, 20.6163, 20.6598, 20.7056, 20.7167, 20.6989, 20.6728, 20.7671, 20.7806, 20.7094, 20.8345, 20.8372, 20.8224, 20.7956, 20.7662, 20.7737, 20.6772, 20.664, 20.6754, 20.7201, 20.6842, 20.5483, 20.5761, 20.5187, 20.4392, 20.5255, 20.5197, 20.5242, 20.5533, 20.5673, 20.5732, 20.5689, 20.6476, 20.631, 20.6102, 20.6005, 20.5914, 20.5843, 20.579, 20.5477, 20.5868, 20.5532, 20.5376, 20.576, 20.6304, 20.6899, 20.7462, 20.7666, 20.7778, 20.7794, 20.695, 20.7085, 20.7281, 20.7166, 20.7353, 20.7674, 20.7722, 20.7708, 20.7574, 20.7379, 20.7269, 20.7383, 20.7623, 20.7657, 20.8034, 20.8056, 20.8038, 20.7903, 20.7993, 20.7971, 20.7993, 20.808, 20.7964, 20.8066, 20.8323, 20.8271, 20.818, 20.8138, 20.8291, 20.8235, 20.8438, 20.841, 20.8909, 20.9641, 20.8477, 20.7513, 20.837, 20.8656, 20.7523, 20.7377, 20.7486, 20.7495, 20.7485, 20.7714, 20.8045, 20.82, 20.7967, 20.7986, 20.8022, 20.82, 20.8263, 20.8481, 20.8796, 20.9604, 20.9632, 20.9834, 20.9747, 20.9336, 20.9548, 20.9443, 20.9656, 20.9358, 20.9468, 20.9564, 20.9622, 20.973, 20.9589, 20.9541, 20.956, 20.9511, 20.963, 20.9534, 20.9423, 20.9586, 20.9639, 20.9637, 20.973, 20.9699, 20.9515, 20.9178, 20.8431, 20.8699, 20.9028, 20.8815, 20.8674, 20.8797, 20.8866, 20.859, 20.8358, 20.8414, 20.851, 20.8637, 20.8472, 20.8577, 20.8671, 20.8687, 20.871, 20.8562, 20.8507, 20.8362, 20.8742, 20.8364, 20.8136, 20.7534, 20.7292, 20.6873, 20.6801, 20.6789, 20.6776, 20.678, 20.6805, 20.6791, 20.685, 20.6878, 20.6883, 20.6901, 20.6917, 20.6909, 20.6911, 20.6932, 20.6919, 20.6943, 20.6937, 20.6967, 20.6967, 20.6958, 20.6975, 20.7013, 20.7003, 20.7021, 20.7, 20.7002, 20.7039, 20.7039, 20.7013, 20.7388, 20.767, 20.8, 20.7505, 20.7289, 20.6998, 20.7226, 20.755, 20.7111, 20.6883, 20.6887, 20.7568, 20.6912, 20.6893, 20.6857, 20.6838, 20.693, 20.6836, 20.7208, 20.7235, 20.6886, 20.6829, 20.6758, 20.7123, 20.6945, 20.8611, 20.7652, 20.898, 20.9165, 20.8788, 20.9223, 20.9334, 20.92, 20.8668, 20.8703, 20.8412, 20.849, 20.8891, 20.9295, 20.8378, 20.8856, 20.8622, 20.8589, 20.8735, 20.8197, 20.8073, 20.85, 20.8538, 20.8174, 20.7768, 20.8268, 20.7079, 20.8247, 20.7706, 20.7576, 20.7852, 20.7369, 20.7105, 20.8252, 20.784, 20.7716, 20.8044, 20.7941, 20.8073, 20.7937, 20.7721, 20.7856, 20.7796, 20.8076, 20.7864, 20.7085, 20.701, 20.735, 20.7393, 20.7647, 20.7405, 20.7224, 20.7028, 20.6948, 20.715, 20.7722, 20.7202, 20.749, 20.7707, 20.7266, 20.7524, 20.7775, 20.7861, 20.7262, 20.7163, 20.7457, 20.7, 20.6542, 20.621, 20.6006, 20.6193, 20.6889, 20.6357, 20.6275, 20.6997, 20.7614, 20.7205, 20.6594, 20.6186, 20.6069, 20.5621, 20.5398, 20.5079, 20.5265, 20.5359, 20.5533, 20.4335, 20.2999, 20.2879, 20.3053, 20.4889, 20.6465, 20.6722, 20.5797, 20.1645, 20.608, 20.6144, 20.5508, 20.6204, 20.7444, 20.6988, 20.651, 20.6608, 20.6896, 20.7196, 20.7013, 20.7289, 20.6435, 20.5843, 20.587, 20.5869, 20.5926, 20.4802, 20.5233, 20.6175, 20.747, 20.749, 20.7484, 20.7639, 20.7209, 20.7024, 20.6765, 20.6526, 20.6694, 20.7391, 20.7561, 20.798, 20.978, 20.979, 20.9816, 20.9982, 20.9964, 20.999, 20.9574, 21.0182, 20.9184, 20.986, 21.0024, 20.9831, 21.0072, 21.0084, 21.0045, 20.9866, 20.9873, 20.9846, 20.9827, 20.9735, 20.9661, 20.9639, 20.9559, 20.9504, 20.9444, 20.9442, 20.9398, 20.9365, 20.932, 20.9284, 20.9262, 20.9235, 20.9083, 20.9111, 20.9086, 20.9025, 20.9042, 20.8888, 20.8784, 20.8783, 20.8607, 20.8785, 20.8785, 20.8447, 20.8634, 20.8366, 20.8582, 20.8328, 20.8362, 20.8258, 20.8415, 20.7769, 20.8232, 20.8308, 20.8299, 20.8472, 20.8608, 20.8481, 20.8427, 20.8542, 20.8547, 20.8582, 20.8553, 20.8509, 20.8581, 20.8482, 20.8343, 20.8154, 20.818, 20.8194, 20.8289, 20.7928, 20.8107, 20.8404, 20.8349, 20.8361, 20.8155, 20.8106, 20.8311, 20.8192, 20.7956, 20.8275, 20.8118, 20.7799, 20.807, 20.7646, 20.6603, 20.5451, 20.644, 20.7449, 20.7903, 20.7791, 20.7526, 20.7483, 20.6681, 20.7349, 20.7681, 20.7948, 20.7246, 20.4395, 20.4338, 20.5408, 20.6102, 20.6038, 20.7042, 20.6904, 20.744, 20.778, 20.7871, 20.7426, 20.557, 20.6944, 20.7043, 20.7317, 20.7075, 20.7663, 20.7257, 20.7158, 20.6287, 20.6585, 20.7174, 20.5976, 20.5846, 20.6285, 20.7557, 20.7694, 20.6284, 20.5973, 20.6855, 20.7007, 20.6721, 20.7585, 20.7476, 20.7229, 20.7249, 20.7076, 20.6675, 20.6672, 20.6848, 20.7148, 20.7667, 20.7629, 20.7773, 20.78, 20.7733, 20.762, 20.7676, 20.7833, 20.8092, 20.8066, 20.8114, 20.8243, 20.8126, 20.7987, 20.7855, 20.7752, 20.7678, 20.7508, 20.7178, 20.666, 20.6768, 20.6517, 20.6442, 20.6534, 20.6617, 20.6664, 20.6714, 20.6595, 20.6807, 20.6922, 20.6861, 20.7005, 20.725, 20.7273, 20.7209, 20.7172, 20.7244, 20.7161, 20.7403, 20.7586, 20.7771, 20.7867, 20.7969, 20.8032, 20.7906, 20.7846, 20.7834, 20.7778, 20.7709, 20.7595, 20.7475, 20.7508, 20.7334, 20.7432, 20.7908, 20.7252, 20.7377, 20.7284, 20.7878, 20.7798, 20.8166, 20.739, 20.687, 20.5466, 20.5461, 20.6069, 20.6241, 20.608, 20.6599, 20.619, 20.5744, 20.4819, 20.4388, 20.4168, 20.4284, 20.4668, 20.4713, 20.5257, 20.4397, 20.4005, 20.4207, 20.4055, 20.4173, 20.4292, 20.5359, 20.4969, 20.5227, 20.487, 20.4624, 20.494, 20.5706, 20.5653, 20.5459, 20.633, 20.7199, 20.6714, 20.7361, 20.7805, 20.7751, 20.7708, 20.7896, 20.8025, 20.7969, 20.7974, 20.8011, 20.8063, 20.813, 20.8121, 20.8125, 20.8105, 20.8066, 20.7992, 20.7583, 20.7856, 20.7754, 20.806, 20.8031, 20.7961, 20.8098, 20.8027, 20.799, 20.7969, 20.7933, 20.8261, 20.8123, 20.8252, 20.8184, 20.818, 20.8167, 20.8192, 20.8162, 20.8, 20.796, 20.8069, 20.8154, 20.8192, 20.8328, 20.8304, 20.838, 20.8529, 20.8572, 20.8603, 20.8643, 20.8659, 20.8727, 20.8727, 20.8597, 20.8631, 20.8688, 20.8775, 20.88, 20.8826, 20.8839, 20.8862, 20.8769, 20.8886, 20.8927, 20.9043, 20.8884, 20.8709, 20.8681, 20.863, 20.8603, 20.8601, 20.8604, 20.8645, 20.8687, 20.8704, 20.8712, 20.8704, 20.8755, 20.8766, 20.877, 20.8736, 20.8594, 20.8619, 20.864, 20.8667, 20.8673, 20.8682, 20.8626, 20.8611, 20.8609, 20.8624, 20.8626, 20.861, 20.8599, 20.8589, 20.8593, 20.8582, 20.8683, 20.8684, 20.8582, 20.8427, 20.8546, 20.8485, 20.8537, 20.8535, 20.8659, 20.8653, 20.8449, 20.8455, 20.8338, 20.8376, 20.8384, 20.8392, 20.8343, 20.8327, 20.809, 20.8006, 20.8439, 20.8377, 20.8355, 20.8402, 20.8492, 20.8682, 20.8629, 20.8491, 20.8303, 20.8025, 20.7029, 20.6338, 20.6797, 20.6709, 20.6915, 20.6702, 20.6732, 20.6182, 20.6017, 20.621, 20.6391, 20.6583, 20.6635, 20.6839, 20.7019, 20.7047, 20.717, 20.7437, 20.7669, 20.7758, 20.8039, 20.817, 20.8343, 20.8541, 20.85, 20.8068, 20.8118, 20.7968, 20.8232, 20.8451, 20.8577, 20.8449, 20.8441, 20.8361, 20.8585, 20.7383, 20.832, 20.7935, 20.7362, 20.8316, 20.8611, 20.8394, 20.8698, 20.8898, 20.8369, 20.8222, 20.7895, 20.7961, 20.8002, 20.7816, 20.8157, 20.705, 20.7199, 20.7724, 20.7029, 20.7912, 20.613, 20.581, 20.7746, 20.7373, 20.7657, 20.7513, 20.4805, 20.5755, 20.7369, 20.6524, 20.6423, 20.7047, 20.6421, 20.7351, 20.7888, 20.759, 20.8261, 20.804, 20.7889, 20.8013, 20.8286, 20.816, 20.76, 20.7476, 20.7446, 20.7095, 20.782, 20.7937, 20.7379, 20.7193, 20.7286, 20.5106, 20.6115, 20.7519, 20.7765, 20.7876, 20.8011, 20.8049, 20.7885, 20.6838, 20.7424, 20.7823, 20.7992, 20.8192, 20.812, 20.838, 20.828, 20.7737, 20.575, 20.444, 20.4226, 20.412, 20.6473, 20.614, 20.7297, 20.7491, 20.7557, 20.7845, 20.7647, 20.7601, 20.7637, 20.7546, 20.6824, 20.7383, 20.7289, 20.7104, 20.6523, 20.6726, 20.7012, 20.6878, 20.7126, 20.5943, 20.4123, 20.6873, 20.7056, 20.6929, 20.6512, 20.6977, 20.5539, 20.6965, 20.715, 20.6519, 20.6772, 20.7172, 20.6549, 20.6371, 20.6823, 20.7421, 20.7108, 20.6469, 20.5919, 20.6164, 20.7195, 20.705, 20.7684, 20.716, 20.6511, 20.6812, 20.6877, 20.7786, 20.7161, 20.6621, 20.7602, 20.8195, 21.0492, 21.01, 21.181, 20.957, 20.7594, 20.69, 20.7739, 20.7412, 21.0373, 20.6513, 21.1429, 21.045, 22.6047, 23.278, 23.549, 23.9744, 23.2331, 22.7068, 22.6621, 22.3843, 22.0349, 21.8274, 21.9826, 22.0103, 22.0559, 22.1042, 22.1804, 22.8156, 24.5968, 25.8325, 25.7912, 25.6392, 27.5845, 27.902, 27.9253, 27.3047, 27.6649, 27.698, 27.6758, 27.639, 27.5939, 27.5362, 27.476, 27.4132, 27.3413, 27.2686, 27.1926, 27.1128, 27.0392, 26.9716, 26.903, 26.8292, 26.7599, 26.6833, 26.6086, 26.5359, 26.4653, 26.4014, 26.3326, 26.2668, 26.1938, 26.1204, 26.0507, 25.9782, 25.904, 25.8265, 25.7466, 25.6648, 25.5812, 25.5002, 25.4223, 25.3485, 25.2705, 25.1964, 25.1251, 25.0555, 24.9891, 24.9238, 24.8578, 24.7964, 24.736, 24.6776, 24.6211, 24.562, 24.5075, 24.4493, 24.3944, 24.3383, 24.2762, 24.2119, 24.145, 24.075, 24.0019, 23.9223, 23.848, 23.7769, 23.7082, 23.6509, 23.5969, 23.5503, 23.5077, 23.4619, 23.4217, 23.3789, 23.3283, 23.2729, 23.2172, 23.1612, 23.1044, 23.0482, 22.9932, 22.9319, 22.8765, 22.8164, 22.7549, 22.6976, 22.6393, 22.5805, 22.5244, 22.4666, 22.4118, 22.358, 22.303, 22.248, 22.1887, 22.1333, 22.0793, 22.0232, 21.9672, 21.9167, 21.8661, 21.8211, 21.7751, 21.732, 21.6918, 21.654, 21.618, 21.583, 21.5497, 21.5199, 21.4918, 21.464, 21.434, 21.4112, 21.3876, 21.3637, 21.351, 21.3424, 21.3363, 21.3328, 21.33, 21.3272, 21.3324, 21.3403, 21.3513, 21.3727, 21.3765, 21.3839, 21.4099, 21.4117, 21.4207, 21.4362, 21.4883, 21.6362, 23.7365, 22.5885, 22.1374, 21.7097, 21.8551, 22.2231, 22.6074, 22.9524, 23.3036, 23.636, 25.9662, 26.2943, 26.5729, 26.7087, 26.7165, 26.7217, 26.6546, 26.607, 26.4167, 25.9872, 25.6544, 25.4122, 25.2069, 25.056, 24.9151, 24.8024, 24.6995, 24.612, 24.5428, 24.4824, 24.4472, 24.4444, 24.4517, 24.4629, 24.4767, 24.4926, 24.509, 24.522, 24.5348, 24.5474, 24.5573, 24.5677, 24.577, 24.5844, 24.5916, 24.5977, 24.6025, 24.6073, 24.6122, 24.6164, 24.6209, 24.6247, 24.6285, 24.6319, 24.6356, 24.6384, 24.6422, 24.6455, 24.6486, 24.6508, 24.6547, 24.6569, 24.6606, 24.6642, 24.6668, 24.6696, 24.6729, 24.6757, 24.6779, 24.6808, 24.6833, 24.6845, 24.6859, 24.6889, 24.6906, 24.6925, 24.6943, 24.6949, 24.6966, 24.6976, 24.6972, 24.6994, 24.6994, 24.7007, 24.7011, 24.7014, 24.7019, 24.7038, 24.7043, 24.705, 24.7047, 24.7068, 24.7062, 24.7065, 24.7076, 24.7078, 24.7079, 24.7097, 24.7098, 24.7106, 24.7087, 24.7089, 24.7107, 24.6519, 24.6079, 24.5706, 24.5327, 24.489, 24.4494, 24.4222, 24.4029, 24.3866, 24.3661, 24.3406, 24.3203, 24.3065, 24.3007, 24.2971, 24.2944, 24.2697, 24.2545, 24.2388, 24.2232, 24.2105, 24.1978, 24.1951, 24.1883, 24.1773, 24.1704, 24.1665, 24.1588, 24.1595, 24.1637, 24.1613, 24.1651, 24.161, 24.1554}
TEMP_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES_REL =
  {35.347, 35.02, 35.29, 35.003, 35.11, 35.453, 35.069, 35.331, 35.192, 34.979, 35.134, 34.979, 35.003, 34.93, 35.372, 35.036, 35.085, 35.363, 35.552, 35.314, 35.412, 35.314, 35.306, 35.306, 35.273, 35.183, 35.126, 35.331, 35.478, 35.249, 35.053, 35.069, 35.527, 35.658, 35.159, 35.388, 35.339, 35.519, 35.445, 35.388, 35.249, 35.167, 35.306, 35.224, 35.404, 35.339, 35.29, 35.437, 35.502, 35.65, 35.314, 35.257, 35.56, 35.699, 35.502, 35.453, 35.29, 35.38, 35.56, 35.306, 35.363, 35.404, 35.552, 35.38, 35.257, 35.323, 35.576, 35.56, 35.388, 35.396, 35.462, 35.642, 35.519, 35.552, 35.625, 35.241, 35.273, 35.543, 35.568, 35.208, 35.535, 35.38, 35.208, 35.543, 35.404, 35.412, 35.282, 35.314, 35.625, 35.29, 35.363, 35.249, 35.552, 35.323, 35.38, 35.339, 35.257, 35.265, 35.282, 35.543, 35.347, 35.093, 35.118, 35.224, 35.543, 35.462, 35.077, 35.208, 35.069, 35.339, 35.126, 35.265, 35.167, 35.421, 35.102, 35.568, 35.249, 35.257, 34.979, 35.012, 34.93, 34.897, 35.167, 35.069, 35.053, 34.979, 34.987, 34.995, 35.053, 34.971, 35.257, 34.881, 34.93, 35.044, 35.151, 35.126, 35.003, 35.151, 34.815, 34.84, 34.93, 35.003, 34.807, 35.167, 34.971, 34.791, 34.954, 35.053, 34.922, 35.265, 35.126, 34.791, 35.085, 35.249, 35.11, 34.979, 34.963, 35.053, 35.183, 35.118, 35.11, 35.069, 35.11, 35.102, 35.306, 35.044, 35.11, 35.2, 35.339, 35.167, 35.159, 35.093, 35.012, 35.126, 35.175, 35.192, 35.265, 35.282, 35.036, 35.282, 35.2, 35.347, 35.233, 35.2, 35.306, 35.421, 35.519, 35.38, 35.241, 35.298, 34.971, 35.355, 35.453, 35.445, 35.273, 35.331, 35.249, 35.347, 35.331, 35.404, 35.38, 35.151, 35.118, 35.445, 35.38, 35.314, 35.249, 35.535, 35.363, 35.396, 35.355, 35.355, 35.061, 35.462, 35.552, 35.617, 35.143, 35.478, 35.192, 35.568, 35.363, 35.216, 35.208, 35.445, 35.282, 35.167, 35.003, 35.192, 35.208, 35.216, 35.355, 35.208, 35.355, 35.126, 35.085, 35.282, 35.453, 35.306, 35.053, 35.249, 35.462, 35.053, 34.873, 35.65, 35.11, 35.143, 35.102, 35.175, 35.053, 35.29, 35.053, 35.012, 35.02, 35.233, 35.012, 34.946, 34.881, 34.987, 35.036, 35.241, 35.028, 35.102, 34.807, 34.824, 34.799, 34.889, 35.175, 34.734, 34.873, 35.02, 34.815, 35.093, 34.652, 35.175, 34.848, 35.159, 34.807, 35.224, 34.799, 35.003, 35.102, 35.175, 34.815, 35.061, 35.012, 34.873, 34.815, 35.003, 34.979, 34.995, 34.774, 34.758, 35.306, 35.093, 35.159, 35.069, 35.257, 34.873, 35.273, 35.077, 35.003, 35.151, 35.134, 35.102, 35.2, 35.257, 35.151, 35.085, 35.167, 35.339, 35.036, 34.897, 35.061, 35.044, 35.061, 35.233, 35.298, 35.331, 35.11, 35.527, 35.224, 34.922, 35.249, 35.208, 35.183, 35.314, 35.453, 35.093, 35.331, 35.306, 35.118, 35.249, 35.372, 35.462, 35.748, 35.282, 35.331, 35.363, 35.404, 35.462, 35.249, 35.47, 35.535, 35.584, 35.421, 35.568, 35.519, 35.429, 35.363, 35.519, 35.421, 35.38, 35.306, 35.421, 35.511, 35.535, 35.527, 35.576, 35.323, 35.642, 35.429, 35.363, 35.306, 35.511, 35.502, 35.821, 35.601, 35.429, 35.396, 35.445, 35.609, 35.92, 35.233, 35.666, 35.854, 35.249, 35.282, 35.265, 35.478, 35.265, 35.437, 35.625, 35.159, 35.208, 35.412, 35.257, 35.167, 35.11, 35.527, 34.954, 35.159, 35.061, 35.511, 35.175, 35.085, 35.462, 35.02, 34.856, 35.151, 35.093, 35.053, 35.233, 35.429, 34.979, 34.922, 34.995, 34.881, 34.946, 34.905, 35.192, 34.824, 34.725, 34.742, 35.143, 34.783, 34.701, 34.971, 35.053, 34.971, 34.954, 34.783, 34.873, 35.126, 35.028, 35.003, 34.611, 34.783, 34.545, 34.963, 34.963, 34.57, 34.742, 34.954, 34.84, 34.799, 34.946, 34.742, 35.077, 35.044, 34.979, 35.249, 34.848, 35.118, 35.29, 34.774, 35.028, 35.044, 34.938, 35.061, 35.404, 35.257, 35.249, 35.134, 35.012, 35.421, 34.979, 34.938, 34.979, 35.183, 34.848, 34.668, 35.388, 35.11, 34.913, 35.314, 34.905, 35.224, 35.372, 35.159, 35.331, 35.527, 35.233, 35.257, 35.183, 35.494, 35.47, 35.363, 35.617, 35.568, 35.682, 35.707, 35.183, 35.306, 35.29, 35.437, 35.306, 35.552, 35.486, 35.486, 35.969, 35.298, 35.494, 35.462, 35.363, 35.527, 35.535, 35.314, 35.805, 35.584, 35.429, 35.306, 35.952, 35.658, 35.388, 35.821, 35.633, 35.511, 35.854, 35.821, 35.494, 35.502, 35.47, 35.216, 35.756, 35.609, 35.592, 35.895, 35.781, 35.707, 35.592, 35.462, 35.601, 35.47, 35.339, 35.216, 35.437, 35.077, 35.445, 35.323, 35.38, 35.462, 35.347, 34.954, 35.061, 34.873, 35.151, 35.453, 35.003, 34.938, 35.134, 35.069, 35.11, 35.134, 35.183, 34.848, 34.873, 35.061, 34.881, 34.676, 34.701, 35.192, 34.873, 34.848, 34.987, 34.39, 34.815, 34.807, 35.028, 35.085, 35.102, 34.684, 34.913, 35.012, 34.954, 35.134, 34.619, 35.085, 34.889, 35.143, 35.003, 35.249, 34.734, 34.824, 35.061, 35.183, 35.044, 35.028, 35.372, 34.979, 34.979, 35.159, 34.717, 35.159, 34.725, 35.02, 35.02, 35.134, 34.905, 35.093, 35.241, 35.478, 35.093, 35.044, 35.331, 35.355, 34.946, 35.552, 35.233, 35.224, 35.306, 34.946, 34.995, 35.126, 35.568, 35.192, 35.012, 35.069, 35.494, 35.249, 35.306, 35.29, 34.987, 35.282, 35.404, 35.813, 35.47, 35.478, 35.609, 35.478, 35.658, 35.535, 35.74, 35.47, 35.2, 35.363, 35.429, 35.486, 35.568, 35.265, 35.388, 35.658, 35.486, 35.102, 35.502, 35.003, 35.543, 35.249, 35.453, 35.314, 35.592, 35.437, 35.462, 35.257, 35.396, 35.543, 35.707, 35.633, 35.453, 35.674, 35.372, 35.83, 35.772, 35.797, 35.568, 35.265, 35.396, 35.355, 35.601, 35.699, 35.478, 35.625, 35.339, 35.462, 35.781, 35.592, 35.601, 35.421, 35.421, 35.323, 35.486, 35.601, 35.028, 35.192, 35.216, 35.175, 35.355, 35.502, 35.282, 35.265, 34.987, 35.134, 35.306, 35.224, 35.257, 35.102, 35.012, 35.069, 35.224, 34.913, 34.954, 35.053, 35.167, 34.783, 35.175, 35.118, 34.75, 34.668, 34.856, 34.709, 35.126, 34.93, 34.979, 34.815, 34.856, 35.069, 34.905, 34.701, 34.791, 35.102, 34.701, 34.873, 34.717, 34.922, 34.913, 34.995, 34.84, 34.881, 34.856, 34.881, 34.766, 34.971, 34.963, 34.815, 34.774, 34.979, 35.38, 34.963, 35.265, 35.102, 35.003, 35.053, 35.38, 35.208, 35.282, 34.889, 35.134, 35.233, 34.971, 35.093, 35.355, 35.388, 35.421, 35.257, 34.946, 35.339, 35.249, 35.061, 35.085, 35.044, 35.38, 35.282, 35.323, 35.012, 35.192, 35.306, 35.323, 35.224, 35.102, 35.11, 35.159, 35.2, 35.143, 35.192, 35.224, 35.339, 35.429, 35.249, 35.404, 35.453, 35.192, 35.249, 35.257, 35.552, 35.061, 35.372, 35.486, 35.355, 35.265, 35.47, 35.494, 35.429, 35.494, 35.478, 35.396, 35.494, 35.584, 35.339, 35.732, 35.38, 35.584, 35.584, 35.543, 35.429, 35.56, 35.601, 35.568, 35.723, 35.527, 35.642, 35.699, 35.666, 35.494, 35.83, 35.609, 35.674, 35.486, 35.781, 35.666, 35.879, 35.699, 35.691, 35.715, 35.797, 35.666, 35.691, 35.666, 35.56, 35.617, 35.74, 35.552, 35.543, 35.47, 35.502, 35.355, 35.568, 35.56, 35.339, 35.396, 35.282, 35.355, 35.216, 35.192, 35.339, 34.987, 35.257, 35.183, 35.257, 35.102, 35.053, 35.167, 35.036, 34.913, 34.954, 35.093, 34.995, 35.159, 35.012, 35.012, 35.028, 35.134, 34.971, 34.897, 34.799, 34.758, 34.791, 34.922, 34.889, 34.979, 34.913, 35.241, 35.003, 35.102, 35.126, 34.963, 35.036, 35.396, 35.118, 35.298, 35.216, 35.061, 35.388, 35.462, 35.183, 35.445, 35.233, 35.273, 35.2, 35.486, 35.502, 35.421, 35.65, 35.633, 35.388, 35.748, 35.633, 35.658, 35.478, 0.516, -0.253, -0.229, -0.237, -0.253, -0.261, -0.261, -0.261, -0.261, -0.261, -0.261, -0.27, -0.261, -0.261, -0.27, -0.261, -0.261, -0.261, -0.261, -0.286, 0.009, 0.0, -0.008, -0.278, -0.032, -0.041, -0.041, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.057, -0.057, -0.057, -0.049, -0.057, -0.057, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.049, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.032, -0.032, -0.041, -0.032, -0.041, -0.032, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.041, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.032, -0.024, -0.032, -0.032, -0.024, -0.024, -0.024, -0.024, -0.024, -0.016, -0.024, -0.024, -0.024, -0.024, -0.024, -0.024, -0.016, -0.016, -0.024, -0.024, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, -0.016, 0.0, -0.245, -0.229, -0.253, -0.253, -0.253, -0.253, -0.261, -0.261, -0.27, -0.253, -0.261, -0.245, -0.253, -0.261, -0.237, -0.245, -0.237, -0.245, -0.237, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.245, -0.237, -0.237, -0.245, -0.237, -0.237, -0.237, -0.237, -0.237, -0.229, -0.229, -0.229, -0.229, -0.229, -0.229, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.229, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.221, -0.229, -0.221, -0.229, -0.229, -0.237, -0.237, -0.221, -0.229, -0.229, -0.229, -0.237, -0.237, -0.237, -0.237, -0.237, -0.237, -0.237, -0.237, -0.245, -0.237, -0.237, -0.237, -0.245, -0.253, -0.245, -0.237, -0.245, -0.245, -0.237, -0.237, -0.229, -0.229, -0.229, -0.237, -0.229, -0.229, -0.229, -0.229, -0.229, -0.229, -0.221, -0.221, -0.229, -0.221, -0.221, -0.221, -0.212, -0.221, -0.221, -0.212, -0.204, -0.212, -0.204, -0.204, -0.204, -0.204, -0.204, -0.204, -0.204, -0.196, -0.196, -0.196, -0.204, -0.204, -0.204, -0.204, -0.204, -0.204, -0.204, -0.212}
PRES_REL_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {35.0965, 34.769646, 35.04206, 34.75952, 34.861603, 35.202053, 34.820747, 35.082924, 34.943333, 34.73225, 34.885437, 34.73225, 34.75952, 34.68804, 35.123764, 34.79013, 34.841232, 35.116993, 35.29731, 35.065884, 35.161198, 35.065884, 35.055656, 35.055656, 35.025036, 34.936546, 34.88209, 35.082924, 35.229317, 35.001198, 34.807156, 34.820747, 35.27695, 35.40974, 34.91271, 35.137363, 35.093155, 35.266712, 35.198708, 35.137363, 35.001198, 34.92295, 35.055656, 34.97394, 35.157852, 35.093155, 35.04206, 35.18846, 35.249695, 35.39949, 35.065884, 35.00455, 35.307556, 35.450592, 35.249695, 35.202053, 35.04206, 35.134018, 35.307556, 35.055656, 35.116993, 35.157852, 35.29731, 35.134018, 35.00455, 35.07267, 35.328033, 35.307556, 35.137363, 35.147602, 35.21572, 35.38925, 35.266712, 35.29731, 35.37223, 34.99441, 35.025036, 35.29054, 35.317802, 34.96381, 35.287193, 35.134018, 34.96381, 35.29054, 35.157852, 35.161198, 35.031815, 35.065884, 35.37223, 35.04206, 35.116993, 35.001198, 35.29731, 35.07267, 35.134018, 35.093155, 35.00455, 35.01479, 35.031815, 35.29054, 35.0965, 34.84459, 34.871853, 34.97394, 35.29054, 35.21572, 34.830994, 34.96381, 34.820747, 35.093155, 34.88209, 35.01479, 34.92295, 35.174877, 34.851364, 35.317802, 35.001198, 35.00455, 34.73225, 34.766304, 34.68804, 34.65053, 34.92295, 34.820747, 34.807156, 34.73225, 34.73903, 34.749275, 34.807156, 34.728905, 35.00455, 34.636948, 34.68804, 34.800385, 34.902462, 34.88209, 34.75952, 34.902462, 34.568813, 34.596073, 34.68804, 34.75952, 34.56547, 34.92295, 34.728905, 34.544964, 34.70842, 34.807156, 34.677803, 35.01479, 34.88209, 34.544964, 34.841232, 35.001198, 34.861603, 34.73225, 34.71866, 34.807156, 34.936546, 34.871853, 34.861603, 34.820747, 34.861603, 34.851364, 35.055656, 34.800385, 34.861603, 34.95357, 35.093155, 34.92295, 34.91271, 34.84459, 34.766304, 34.88209, 34.9263, 34.943333, 35.01479, 35.031815, 34.79013, 35.031815, 34.95357, 35.0965, 34.984173, 34.95357, 35.055656, 35.174877, 35.266712, 35.134018, 34.99441, 35.052307, 34.728905, 35.106747, 35.202053, 35.198708, 35.025036, 35.082924, 35.001198, 35.0965, 35.082924, 35.157852, 35.134018, 34.902462, 34.871853, 35.198708, 35.134018, 35.065884, 35.001198, 35.287193, 35.116993, 35.147602, 35.106747, 35.106747, 34.810493, 35.21572, 35.29731, 35.36889, 34.899113, 35.229317, 34.943333, 35.317802, 35.116993, 34.967148, 34.96381, 35.198708, 35.031815, 34.92295, 34.75952, 34.943333, 34.96381, 34.967148, 35.106747, 34.96381, 35.106747, 34.88209, 34.841232, 35.031815, 35.202053, 35.055656, 34.807156, 35.001198, 35.21572, 34.807156, 34.626694, 35.39949, 34.861603, 34.899113, 34.851364, 34.9263, 34.807156, 35.04206, 34.807156, 34.766304, 34.769646, 34.984173, 34.766304, 34.70164, 34.636948, 34.73903, 34.79013, 34.99441, 34.779892, 34.851364, 34.56547, 34.57558, 34.55521, 34.647186, 34.9263, 34.49397, 34.626694, 34.769646, 34.568813, 34.84459, 34.41225, 34.9263, 34.606323, 34.91271, 34.56547, 34.97394, 34.55521, 34.75952, 34.851364, 34.9263, 34.568813, 34.810493, 34.766304, 34.626694, 34.568813, 34.75952, 34.73225, 34.749275, 34.52795, 34.514366, 35.055656, 34.84459, 34.91271, 34.820747, 35.00455, 34.626694, 35.025036, 34.830994, 34.75952, 34.902462, 34.885437, 34.851364, 34.95357, 35.00455, 34.902462, 34.841232, 34.92295, 35.093155, 34.79013, 34.65053, 34.810493, 34.800385, 34.810493, 34.984173, 35.052307, 35.082924, 34.861603, 35.27695, 34.97394, 34.677803, 35.001198, 34.96381, 34.936546, 35.065884, 35.202053, 34.84459, 35.082924, 35.055656, 34.871853, 35.001198, 35.123764, 35.21572, 35.49479, 35.031815, 35.082924, 35.116993, 35.157852, 35.21572, 35.001198, 35.21907, 35.287193, 35.331383, 35.174877, 35.317802, 35.266712, 35.178223, 35.116993, 35.266712, 35.174877, 35.134018, 35.055656, 35.174877, 35.259926, 35.287193, 35.27695, 35.328033, 35.07267, 35.38925, 35.178223, 35.116993, 35.055656, 35.259926, 35.249695, 35.56626, 35.348396, 35.178223, 35.147602, 35.198708, 35.358643, 35.66498, 34.984173, 35.413086, 35.603756, 35.001198, 35.031815, 35.01479, 35.229317, 35.01479, 35.18846, 35.37223, 34.91271, 34.96381, 35.161198, 35.00455, 34.92295, 34.861603, 35.27695, 34.70842, 34.91271, 34.810493, 35.259926, 34.9263, 34.841232, 35.21572, 34.769646, 34.609676, 34.902462, 34.84459, 34.807156, 34.984173, 35.178223, 34.73225, 34.677803, 34.749275, 34.636948, 34.70164, 34.66077, 34.943333, 34.57558, 34.476837, 34.497326, 34.899113, 34.534725, 34.456474, 34.728905, 34.807156, 34.728905, 34.70842, 34.534725, 34.626694, 34.88209, 34.779892, 34.75952, 34.3645, 34.534725, 34.303265, 34.71866, 34.71866, 34.323643, 34.497326, 34.70842, 34.596073, 34.55521, 34.70164, 34.497326, 34.830994, 34.800385, 34.73225, 35.001198, 34.606323, 34.871853, 35.04206, 34.52795, 34.779892, 34.800385, 34.691387, 34.810493, 35.157852, 35.00455, 35.001198, 34.885437, 34.766304, 35.174877, 34.73225, 34.691387, 34.73225, 34.936546, 34.606323, 34.42585, 35.137363, 34.861603, 34.671017, 35.065884, 34.66077, 34.97394, 35.123764, 34.91271, 35.082924, 35.27695, 34.984173, 35.00455, 34.936546, 35.246346, 35.21907, 35.116993, 35.36889, 35.317802, 35.433567, 35.45394, 34.936546, 35.055656, 35.04206, 35.18846, 35.055656, 35.29731, 35.239555, 35.239555, 35.716064, 35.052307, 35.246346, 35.21572, 35.116993, 35.27695, 35.287193, 35.065884, 35.552677, 35.331383, 35.178223, 35.055656, 35.699055, 35.40974, 35.137363, 35.56626, 35.382477, 35.259926, 35.603756, 35.56626, 35.246346, 35.249695, 35.21907, 34.967148, 35.501568, 35.358643, 35.341625, 35.64461, 35.532307, 35.45394, 35.341625, 35.21572, 35.348396, 35.21907, 35.093155, 34.967148, 35.18846, 34.830994, 35.198708, 35.07267, 35.134018, 35.21572, 35.0965, 34.70842, 34.810493, 34.626694, 34.902462, 35.202053, 34.75952, 34.691387, 34.885437, 34.820747, 34.861603, 34.885437, 34.936546, 34.606323, 34.626694, 34.810493, 34.636948, 34.436096, 34.456474, 34.943333, 34.626694, 34.606323, 34.73903, 34.150055, 34.568813, 34.56547, 34.779892, 34.841232, 34.851364, 34.435974, 34.671017, 34.766304, 34.70842, 34.885437, 34.374752, 34.841232, 34.647186, 34.899113, 34.75952, 35.001198, 34.49397, 34.57558, 34.810493, 34.936546, 34.800385, 34.779892, 35.123764, 34.73225, 34.73225, 34.91271, 34.47349, 34.91271, 34.476837, 34.769646, 34.769646, 34.885437, 34.66077, 34.84459, 34.99441, 35.229317, 34.84459, 34.800385, 35.082924, 35.106747, 34.70164, 35.29731, 34.984173, 34.97394, 35.055656, 34.70164, 34.749275, 34.88209, 35.317802, 34.943333, 34.766304, 34.820747, 35.246346, 35.001198, 35.055656, 35.04206, 34.73903, 35.031815, 35.157852, 35.562916, 35.21907, 35.229317, 35.358643, 35.229317, 35.40974, 35.287193, 35.491447, 35.21907, 34.95357, 35.116993, 35.178223, 35.239555, 35.317802, 35.01479, 35.137363, 35.40974, 35.239555, 34.851364, 35.249695, 34.75952, 35.29054, 35.001198, 35.202053, 35.065884, 35.341625, 35.18846, 35.21572, 35.00455, 35.147602, 35.29054, 35.45394, 35.382477, 35.202053, 35.42333, 35.123764, 35.579933, 35.522057, 35.542427, 35.317802, 35.01479, 35.147602, 35.106747, 35.348396, 35.450592, 35.229317, 35.37223, 35.093155, 35.21572, 35.532307, 35.341625, 35.348396, 35.174877, 35.174877, 35.07267, 35.239555, 35.348396, 34.779892, 34.943333, 34.967148, 34.9263, 35.106747, 35.249695, 35.031815, 35.01479, 34.73903, 34.885437, 35.055656, 34.97394, 35.00455, 34.851364, 34.766304, 34.820747, 34.97394, 34.671017, 34.70842, 34.807156, 34.92295, 34.534725, 34.9263, 34.871853, 34.504116, 34.42585, 34.609676, 34.466717, 34.88209, 34.68804, 34.73225, 34.568813, 34.609676, 34.820747, 34.66077, 34.456474, 34.544964, 34.851364, 34.456474, 34.626694, 34.47349, 34.677803, 34.671017, 34.749275, 34.596073, 34.636948, 34.609676, 34.636948, 34.5177, 34.728905, 34.71866, 34.568813, 34.52795, 34.73225, 35.134018, 34.71866, 35.01479, 34.851364, 34.75952, 34.807156, 35.134018, 34.96381, 35.031815, 34.647186, 34.885437, 34.984173, 34.728905, 34.84459, 35.106747, 35.137363, 35.174877, 35.00455, 34.70164, 35.093155, 35.001198, 34.810493, 34.841232, 34.800385, 35.134018, 35.031815, 35.07267, 34.766304, 34.943333, 35.055656, 35.07267, 34.97394, 34.851364, 34.861603, 34.91271, 34.95357, 34.899113, 34.943333, 34.97394, 35.093155, 35.178223, 35.001198, 35.157852, 35.202053, 34.943333, 35.001198, 35.00455, 35.29731, 34.810493, 35.123764, 35.239555, 35.106747, 35.01479, 35.21907, 35.246346, 35.178223, 35.246346, 35.229317, 35.147602, 35.246346, 35.331383, 35.093155, 35.481194, 35.134018, 35.331383, 35.331383, 35.29054, 35.178223, 35.307556, 35.348396, 35.317802, 35.474426, 35.27695, 35.38925, 35.450592, 35.413086, 35.246346, 35.579933, 35.358643, 35.42333, 35.239555, 35.532307, 35.413086, 35.62412, 35.450592, 35.44035, 35.464188, 35.542427, 35.413086, 35.44035, 35.413086, 35.307556, 35.36889, 35.491447, 35.29731, 35.29054, 35.21907, 35.249695, 35.106747, 35.317802, 35.307556, 35.093155, 35.147602, 35.031815, 35.106747, 34.967148, 34.943333, 35.093155, 34.73903, 35.00455, 34.936546, 35.00455, 34.851364, 34.807156, 34.92295, 34.79013, 34.671017, 34.70842, 34.84459, 34.749275, 34.91271, 34.766304, 34.766304, 34.779892, 34.885437, 34.728905, 34.65053, 34.55521, 34.514366, 34.544964, 34.677803, 34.647186, 34.73225, 34.671017, 34.99441, 34.75952, 34.851364, 34.88209, 34.71866, 34.79013, 35.147602, 34.871853, 35.052307, 34.967148, 34.810493, 35.137363, 35.21572, 34.936546, 35.198708, 34.984173, 35.025036, 34.95357, 35.239555, 35.249695, 35.174877, 35.39949, 35.382477, 35.137363, 35.49479, 35.382477, 35.40974, 35.229317, 0.5152711, -0.24732095, -0.2267286, -0.23705038, -0.24732095, -0.26109928, -0.26109928, -0.26109928, -0.26109928, -0.26109928, -0.26109928, -0.26795742, -0.26109928, -0.26109928, -0.26795742, -0.26109928, -0.26109928, -0.26109928, -0.26109928, -0.285143, 0.0068574273, 0.0, -0.0034065007, -0.27827927, -0.034368884, -0.0412264, -0.0412264, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.058411002, -0.058411002, -0.058411002, -0.044633, -0.058411002, -0.058411002, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.044633, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.034368884, -0.034368884, -0.0412264, -0.034368884, -0.0412264, -0.034368884, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.0412264, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.034368884, -0.020590948, -0.034368884, -0.034368884, -0.020590948, -0.020590948, -0.020590948, -0.020590948, -0.020590948, -0.017184408, -0.020590948, -0.020590948, -0.020590948, -0.020590948, -0.020590948, -0.020590948, -0.017184408, -0.017184408, -0.020590948, -0.020590948, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, -0.017184408, 0.0, -0.24391396, -0.2267286, -0.24732095, -0.24732095, -0.24732095, -0.24732095, -0.26109928, -0.26109928, -0.26795742, -0.24732095, -0.26109928, -0.24391396, -0.24732095, -0.26109928, -0.23705038, -0.24391396, -0.23705038, -0.24391396, -0.23705038, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.24391396, -0.23705038, -0.23705038, -0.24391396, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.2267286, -0.2267286, -0.2267286, -0.2267286, -0.2267286, -0.2267286, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2267286, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2233216, -0.2267286, -0.2233216, -0.2267286, -0.2267286, -0.23705038, -0.23705038, -0.2233216, -0.2267286, -0.2267286, -0.2267286, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.23705038, -0.24391396, -0.23705038, -0.23705038, -0.23705038, -0.24391396, -0.24732095, -0.24391396, -0.23705038, -0.24391396, -0.24391396, -0.23705038, -0.23705038, -0.2267286, -0.2267286, -0.2267286, -0.23705038, -0.2267286, -0.2267286, -0.2267286, -0.2267286, -0.2267286, -0.2267286, -0.2233216, -0.2233216, -0.2267286, -0.2233216, -0.2233216, -0.2233216, -0.21300706, -0.2233216, -0.2233216, -0.21300706, -0.20268539, -0.21300706, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.19582188, -0.19582188, -0.19582188, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.20268539, -0.21300706}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
