netcdf file-165.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (27 currently)
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074, 22530.036261574074}
TEMP =
  {21.9219, 21.9138, 21.8967, 21.8763, 21.8575, 21.8339, 21.8203, 21.8173, 21.8158, 21.8141, 21.8113, 21.8109, 21.8106, 21.8083, 21.8072, 21.8068, 21.8064, 21.8062, 21.8058, 21.8055, 21.8055, 21.8058, 21.806, 21.806, 21.8064, 21.8068, 21.8088}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
