netcdf file-155.nc {
  dimensions:
    DEPTH = 24;
  variables:
    float LATITUDE(DEPTH=24);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=24);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=24);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=24);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=24);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=24);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074, 22166.08699074074}
TEMP =
  {24.5057, 24.5043, 24.4974, 24.4892, 24.4721, 24.4447, 24.4172, 24.3927, 24.3733, 24.3589, 24.35, 24.344, 24.3384, 24.3338, 24.3307, 24.3282, 24.3266, 24.3257, 24.3251, 24.3246, 24.3242, 24.3243, 24.3238, 24.3232}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.854}
}
