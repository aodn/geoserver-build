netcdf file-73.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (46 currently)
  variables:
    float LATITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=46);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=46);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=46);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=46);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875, 22696.0875}
TEMP =
  {23.623356, 23.541893, 23.520237, 23.515057, 23.519209, 23.515104, 23.516766, 23.504606, 23.50376, 23.49967, 23.501575, 23.501358, 23.502605, 23.512085, 23.513294, 23.510876, 23.506853, 23.513098, 23.510168, 23.511484, 23.513588, 23.510727, 23.507465, 23.50685, 23.507761, 23.501036, 23.50052, 23.479483, 23.475851, 23.46883, 23.464346, 23.418505, 23.39537, 23.30084, 22.912512, 22.693594, 22.543201, 22.504702, 22.49081, 22.459059, 22.45267, 22.4592, 22.448185, 22.437868, 22.440351, 22.44105}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0}
}
