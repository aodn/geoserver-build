netcdf IMOS_ANMN-TS_20150113T230000Z_WATR20_FV01_WATR20-1407-RBR-DR1050P-196_END-20150120T071600Z_id-7742.nc {
  dimensions:
    TIME = UNLIMITED;   // (4569 currently)
  variables:
    double TIME(TIME=4569);
      :standard_name = "time";
      :long_name = "time";
      :units = "days since 1950-01-01 00:00:00 UTC";
      :calendar = "gregorian";
      :axis = "T";
      :valid_min = 0.0; // double
      :valid_max = 90000.0; // double

    double LATITUDE;
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees north";
      :axis = "Y";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -90.0; // double
      :valid_max = 90.0; // double

    double LONGITUDE;
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees east";
      :axis = "X";
      :reference_datum = "geographical coordinates, WGS84 projection";
      :valid_min = -180.0; // double
      :valid_max = 180.0; // double

    float NOMINAL_DEPTH;
      :standard_name = "depth";
      :long_name = "nominal depth";
      :units = "metres";
      :axis = "Z";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float

    float TEMP(TIME=4569);
      :standard_name = "sea_water_temperature";
      :long_name = "sea_water_temperature";
      :units = "Celsius";
      :valid_min = -2.5f; // float
      :valid_max = 40.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "TEMP_quality_control";

    byte TEMP_quality_control(TIME=4569);
      :standard_name = "sea_water_temperature status_flag";
      :long_name = "quality flag for sea_water_temperature";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1.0; // double
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float CNDC(TIME=4569);
      :standard_name = "sea_water_electrical_conductivity";
      :long_name = "sea_water_electrical_conductivity";
      :units = "S m-1";
      :valid_min = 0.0f; // float
      :valid_max = 50000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "CNDC_quality_control";

    byte CNDC_quality_control(TIME=4569);
      :standard_name = "sea_water_electrical_conductivity status_flag";
      :long_name = "quality flag for sea_water_electrical_conductivity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PSAL(TIME=4569);
      :standard_name = "sea_water_salinity";
      :long_name = "sea_water_salinity";
      :units = "1e-3";
      :valid_min = 2.0f; // float
      :valid_max = 41.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PSAL_quality_control";

    byte PSAL_quality_control(TIME=4569);
      :standard_name = "sea_water_salinity status_flag";
      :long_name = "quality flag for sea_water_salinity";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES(TIME=4569);
      :standard_name = "sea_water_pressure";
      :long_name = "sea_water_pressure";
      :units = "dbar";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_quality_control";

    byte PRES_quality_control(TIME=4569);
      :standard_name = "sea_water_pressure status_flag";
      :long_name = "quality flag for sea_water_pressure";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float PRES_REL(TIME=4569);
      :standard_name = "sea_water_pressure_due_to_sea_water";
      :long_name = "sea_water_pressure_due_to_sea_water";
      :units = "dbar";
      :valid_min = -15.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE NOMINAL_DEPTH DEPTH";
      :ancillary_variables = "PRES_REL_quality_control";

    byte PRES_REL_quality_control(TIME=4569);
      :standard_name = "sea_water_pressure_due_to_sea_water status_flag";
      :long_name = "quality flag for sea_water_pressure_due_to_sea_water";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

    float DEPTH(TIME=4569);
      :standard_name = "depth";
      :long_name = "depth";
      :units = "metres";
      :positive = "down";
      :reference_datum = "sea surface";
      :valid_min = -5.0f; // float
      :valid_max = 12000.0f; // float
      :_FillValue = 999999.0f; // float
      :ancillary_variables = "DEPTH_quality_control";

    byte DEPTH_quality_control(TIME=4569);
      :standard_name = "depth status_flag";
      :long_name = "quality flag for depth";
      :valid_min = 0B; // byte
      :valid_max = 9B; // byte
      :_FillValue = 99B; // byte
      :quality_control_set = 1; // int
      :quality_control_conventions = "IMOS standard set using the IODE flags";
      :flag_values = 0B, 1B, 2B, 3B, 4B, 5B, 6B, 7B, 8B, 9B; // byte
      :flag_meaning = "No_QC_performed Good_data Probably_good_data Bad_data_that_are_potentially_correctable Bad_data Value_changed Not_used Not_used Not_used Missing_value";

  // global attributes:
  :toolbox_version = "2.3b - PCWIN";
  :file_version = "Level 1 - Quality Controlled Data";
  :file_version_quality_control = "Quality controlled data have passed quality assurance procedures such as automated or visual inspection and removal of obvious errors. The data are using standard SI metric units with calibration and other routine pre-processing applied, all time and location values are in absolute coordinates to agreed to standards and datum, metadata exists for the data or for the higher level dataset that the data belongs to. This is the standard IMOS data level and is what should be made available to eMII and to the IMOS community.";
  :project = "Integrated Marine Observing System (IMOS)";
  :Conventions = "CF-1.6,IMOS-1.3";
  :standard_name_vocabulary = "CF-1.6";
  :comment = "Geospatial vertical min/max information has been computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and absolute pressure measurements to which a nominal value for atmospheric pressure (10.1325 dbar) has been substracted.";
  :instrument = "RBR DR1050P";
  :references = "http://www.imos.org.au";
  :site_code = "WATR20";
  :platform_code = "WATR20";
  :deployment_code = "WATR20-1407";
  :featureType = "timeSeries";
  :naming_authority = "IMOS";
  :instrument_serial_number = "14551";
  :history = "2015-01-29T06:31:59Z - depthPP: Depth computed using the Gibbs-SeaWater toolbox (TEOS-10) v3.02 from latitude and absolute pressure measurements to which a nominal value for atmospheric pressure (10.1325 dbar) has been substracted.";
  :geospatial_lat_min = -31.7285666667; // double
  :geospatial_lat_max = -31.7285666667; // double
  :geospatial_lon_min = 115.0371; // double
  :geospatial_lon_max = 115.0371; // double
  :instrument_nominal_depth = 196.0f; // float
  :site_nominal_depth = 210.0f; // float
  :geospatial_vertical_min = -0.068716735f; // float
  :geospatial_vertical_max = 207.40262f; // float
  :geospatial_vertical_positive = "down";
  :time_deployment_start = "2014-07-10T05:00:00Z";
  :time_deployment_end = "2015-01-20T02:40:00Z";
  :time_coverage_start = "2015-01-13T23:00:00Z";
  :time_coverage_end = "2015-01-20T07:16:00Z";
  :data_centre = "eMarine Information Infrastructure (eMII)";
  :data_centre_email = "info@aodn.org.au";
  :institution_references = "http://www.imos.org.au/emii.html";
  :institution = "The citation in a list of references is: \"IMOS [year-of-data-download], [Title], [data-access-url], accessed [date-of-access]\"";
  :acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and and the Super Science Initiative.\"";
  :distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose.";
  :project_acknowledgement = "The collection of this data was funded by IMOS";
 data:
TIME =
  {23753.958333333332, 23753.959722222222, 23753.96111111111, 23753.9625, 23753.963888888888, 23753.965277777777, 23753.966666666667, 23753.968055555557, 23753.969444444443, 23753.970833333333, 23753.972222222223, 23753.973611111112, 23753.975, 23753.97638888889, 23753.977777777778, 23753.979166666668, 23753.980555555554, 23753.981944444444, 23753.983333333334, 23753.984722222223, 23753.98611111111, 23753.9875, 23753.98888888889, 23753.99027777778, 23753.991666666665, 23753.993055555555, 23753.994444444445, 23753.995833333334, 23753.99722222222, 23753.99861111111, 23754.0, 23754.00138888889, 23754.00277777778, 23754.004166666666, 23754.005555555555, 23754.006944444445, 23754.008333333335, 23754.00972222222, 23754.01111111111, 23754.0125, 23754.01388888889, 23754.015277777777, 23754.016666666666, 23754.018055555556, 23754.019444444446, 23754.020833333332, 23754.022222222222, 23754.02361111111, 23754.025, 23754.026388888888, 23754.027777777777, 23754.029166666667, 23754.030555555557, 23754.031944444443, 23754.033333333333, 23754.034722222223, 23754.036111111112, 23754.0375, 23754.03888888889, 23754.040277777778, 23754.041666666668, 23754.043055555554, 23754.044444444444, 23754.045833333334, 23754.047222222223, 23754.04861111111, 23754.05, 23754.05138888889, 23754.05277777778, 23754.054166666665, 23754.055555555555, 23754.056944444445, 23754.058333333334, 23754.05972222222, 23754.06111111111, 23754.0625, 23754.06388888889, 23754.06527777778, 23754.066666666666, 23754.068055555555, 23754.069444444445, 23754.070833333335, 23754.07222222222, 23754.07361111111, 23754.075, 23754.07638888889, 23754.077777777777, 23754.079166666666, 23754.080555555556, 23754.081944444446, 23754.083333333332, 23754.084722222222, 23754.08611111111, 23754.0875, 23754.088888888888, 23754.090277777777, 23754.091666666667, 23754.093055555557, 23754.094444444443, 23754.095833333333, 23754.097222222223, 23754.098611111112, 23754.1, 23754.10138888889, 23754.102777777778, 23754.104166666668, 23754.105555555554, 23754.106944444444, 23754.108333333334, 23754.109722222223, 23754.11111111111, 23754.1125, 23754.11388888889, 23754.11527777778, 23754.116666666665, 23754.118055555555, 23754.119444444445, 23754.120833333334, 23754.12222222222, 23754.12361111111, 23754.125, 23754.12638888889, 23754.12777777778, 23754.129166666666, 23754.130555555555, 23754.131944444445, 23754.133333333335, 23754.13472222222, 23754.13611111111, 23754.1375, 23754.13888888889, 23754.140277777777, 23754.141666666666, 23754.143055555556, 23754.144444444446, 23754.145833333332, 23754.147222222222, 23754.14861111111, 23754.15, 23754.151388888888, 23754.152777777777, 23754.154166666667, 23754.155555555557, 23754.156944444443, 23754.158333333333, 23754.159722222223, 23754.161111111112, 23754.1625, 23754.16388888889, 23754.165277777778, 23754.166666666668, 23754.168055555554, 23754.169444444444, 23754.170833333334, 23754.172222222223, 23754.17361111111, 23754.175, 23754.17638888889, 23754.17777777778, 23754.179166666665, 23754.180555555555, 23754.181944444445, 23754.183333333334, 23754.18472222222, 23754.18611111111, 23754.1875, 23754.18888888889, 23754.19027777778, 23754.191666666666, 23754.193055555555, 23754.194444444445, 23754.195833333335, 23754.19722222222, 23754.19861111111, 23754.2, 23754.20138888889, 23754.202777777777, 23754.204166666666, 23754.205555555556, 23754.206944444446, 23754.208333333332, 23754.209722222222, 23754.21111111111, 23754.2125, 23754.213888888888, 23754.215277777777, 23754.216666666667, 23754.218055555557, 23754.219444444443, 23754.220833333333, 23754.222222222223, 23754.223611111112, 23754.225, 23754.22638888889, 23754.227777777778, 23754.229166666668, 23754.230555555554, 23754.231944444444, 23754.233333333334, 23754.234722222223, 23754.23611111111, 23754.2375, 23754.23888888889, 23754.24027777778, 23754.241666666665, 23754.243055555555, 23754.244444444445, 23754.245833333334, 23754.24722222222, 23754.24861111111, 23754.25, 23754.25138888889, 23754.25277777778, 23754.254166666666, 23754.255555555555, 23754.256944444445, 23754.258333333335, 23754.25972222222, 23754.26111111111, 23754.2625, 23754.26388888889, 23754.265277777777, 23754.266666666666, 23754.268055555556, 23754.269444444446, 23754.270833333332, 23754.272222222222, 23754.27361111111, 23754.275, 23754.276388888888, 23754.277777777777, 23754.279166666667, 23754.280555555557, 23754.281944444443, 23754.283333333333, 23754.284722222223, 23754.286111111112, 23754.2875, 23754.28888888889, 23754.290277777778, 23754.291666666668, 23754.293055555554, 23754.294444444444, 23754.295833333334, 23754.297222222223, 23754.29861111111, 23754.3, 23754.30138888889, 23754.30277777778, 23754.304166666665, 23754.305555555555, 23754.306944444445, 23754.308333333334, 23754.30972222222, 23754.31111111111, 23754.3125, 23754.31388888889, 23754.31527777778, 23754.316666666666, 23754.318055555555, 23754.319444444445, 23754.320833333335, 23754.32222222222, 23754.32361111111, 23754.325, 23754.32638888889, 23754.327777777777, 23754.329166666666, 23754.330555555556, 23754.331944444446, 23754.333333333332, 23754.334722222222, 23754.33611111111, 23754.3375, 23754.338888888888, 23754.340277777777, 23754.341666666667, 23754.343055555557, 23754.344444444443, 23754.345833333333, 23754.347222222223, 23754.348611111112, 23754.35, 23754.35138888889, 23754.352777777778, 23754.354166666668, 23754.355555555554, 23754.356944444444, 23754.358333333334, 23754.359722222223, 23754.36111111111, 23754.3625, 23754.36388888889, 23754.36527777778, 23754.366666666665, 23754.368055555555, 23754.369444444445, 23754.370833333334, 23754.37222222222, 23754.37361111111, 23754.375, 23754.37638888889, 23754.37777777778, 23754.379166666666, 23754.380555555555, 23754.381944444445, 23754.383333333335, 23754.38472222222, 23754.38611111111, 23754.3875, 23754.38888888889, 23754.390277777777, 23754.391666666666, 23754.393055555556, 23754.394444444446, 23754.395833333332, 23754.397222222222, 23754.39861111111, 23754.4, 23754.401388888888, 23754.402777777777, 23754.404166666667, 23754.405555555557, 23754.406944444443, 23754.408333333333, 23754.409722222223, 23754.411111111112, 23754.4125, 23754.41388888889, 23754.415277777778, 23754.416666666668, 23754.418055555554, 23754.419444444444, 23754.420833333334, 23754.422222222223, 23754.42361111111, 23754.425, 23754.42638888889, 23754.42777777778, 23754.429166666665, 23754.430555555555, 23754.431944444445, 23754.433333333334, 23754.43472222222, 23754.43611111111, 23754.4375, 23754.43888888889, 23754.44027777778, 23754.441666666666, 23754.443055555555, 23754.444444444445, 23754.445833333335, 23754.44722222222, 23754.44861111111, 23754.45, 23754.45138888889, 23754.452777777777, 23754.454166666666, 23754.455555555556, 23754.456944444446, 23754.458333333332, 23754.459722222222, 23754.46111111111, 23754.4625, 23754.463888888888, 23754.465277777777, 23754.466666666667, 23754.468055555557, 23754.469444444443, 23754.470833333333, 23754.472222222223, 23754.473611111112, 23754.475, 23754.47638888889, 23754.477777777778, 23754.479166666668, 23754.480555555554, 23754.481944444444, 23754.483333333334, 23754.484722222223, 23754.48611111111, 23754.4875, 23754.48888888889, 23754.49027777778, 23754.491666666665, 23754.493055555555, 23754.494444444445, 23754.495833333334, 23754.49722222222, 23754.49861111111, 23754.5, 23754.50138888889, 23754.50277777778, 23754.504166666666, 23754.505555555555, 23754.506944444445, 23754.508333333335, 23754.50972222222, 23754.51111111111, 23754.5125, 23754.51388888889, 23754.515277777777, 23754.516666666666, 23754.518055555556, 23754.519444444446, 23754.520833333332, 23754.522222222222, 23754.52361111111, 23754.525, 23754.526388888888, 23754.527777777777, 23754.529166666667, 23754.530555555557, 23754.531944444443, 23754.533333333333, 23754.534722222223, 23754.536111111112, 23754.5375, 23754.53888888889, 23754.540277777778, 23754.541666666668, 23754.543055555554, 23754.544444444444, 23754.545833333334, 23754.547222222223, 23754.54861111111, 23754.55, 23754.55138888889, 23754.55277777778, 23754.554166666665, 23754.555555555555, 23754.556944444445, 23754.558333333334, 23754.55972222222, 23754.56111111111, 23754.5625, 23754.56388888889, 23754.56527777778, 23754.566666666666, 23754.568055555555, 23754.569444444445, 23754.570833333335, 23754.57222222222, 23754.57361111111, 23754.575, 23754.57638888889, 23754.577777777777, 23754.579166666666, 23754.580555555556, 23754.581944444446, 23754.583333333332, 23754.584722222222, 23754.58611111111, 23754.5875, 23754.588888888888, 23754.590277777777, 23754.591666666667, 23754.593055555557, 23754.594444444443, 23754.595833333333, 23754.597222222223, 23754.598611111112, 23754.6, 23754.60138888889, 23754.602777777778, 23754.604166666668, 23754.605555555554, 23754.606944444444, 23754.608333333334, 23754.609722222223, 23754.61111111111, 23754.6125, 23754.61388888889, 23754.61527777778, 23754.616666666665, 23754.618055555555, 23754.619444444445, 23754.620833333334, 23754.62222222222, 23754.62361111111, 23754.625, 23754.62638888889, 23754.62777777778, 23754.629166666666, 23754.630555555555, 23754.631944444445, 23754.633333333335, 23754.63472222222, 23754.63611111111, 23754.6375, 23754.63888888889, 23754.640277777777, 23754.641666666666, 23754.643055555556, 23754.644444444446, 23754.645833333332, 23754.647222222222, 23754.64861111111, 23754.65, 23754.651388888888, 23754.652777777777, 23754.654166666667, 23754.655555555557, 23754.656944444443, 23754.658333333333, 23754.659722222223, 23754.661111111112, 23754.6625, 23754.66388888889, 23754.665277777778, 23754.666666666668, 23754.668055555554, 23754.669444444444, 23754.670833333334, 23754.672222222223, 23754.67361111111, 23754.675, 23754.67638888889, 23754.67777777778, 23754.679166666665, 23754.680555555555, 23754.681944444445, 23754.683333333334, 23754.68472222222, 23754.68611111111, 23754.6875, 23754.68888888889, 23754.69027777778, 23754.691666666666, 23754.693055555555, 23754.694444444445, 23754.695833333335, 23754.69722222222, 23754.69861111111, 23754.7, 23754.70138888889, 23754.702777777777, 23754.704166666666, 23754.705555555556, 23754.706944444446, 23754.708333333332, 23754.709722222222, 23754.71111111111, 23754.7125, 23754.713888888888, 23754.715277777777, 23754.716666666667, 23754.718055555557, 23754.719444444443, 23754.720833333333, 23754.722222222223, 23754.723611111112, 23754.725, 23754.72638888889, 23754.727777777778, 23754.729166666668, 23754.730555555554, 23754.731944444444, 23754.733333333334, 23754.734722222223, 23754.73611111111, 23754.7375, 23754.73888888889, 23754.74027777778, 23754.741666666665, 23754.743055555555, 23754.744444444445, 23754.745833333334, 23754.74722222222, 23754.74861111111, 23754.75, 23754.75138888889, 23754.75277777778, 23754.754166666666, 23754.755555555555, 23754.756944444445, 23754.758333333335, 23754.75972222222, 23754.76111111111, 23754.7625, 23754.76388888889, 23754.765277777777, 23754.766666666666, 23754.768055555556, 23754.769444444446, 23754.770833333332, 23754.772222222222, 23754.77361111111, 23754.775, 23754.776388888888, 23754.777777777777, 23754.779166666667, 23754.780555555557, 23754.781944444443, 23754.783333333333, 23754.784722222223, 23754.786111111112, 23754.7875, 23754.78888888889, 23754.790277777778, 23754.791666666668, 23754.793055555554, 23754.794444444444, 23754.795833333334, 23754.797222222223, 23754.79861111111, 23754.8, 23754.80138888889, 23754.80277777778, 23754.804166666665, 23754.805555555555, 23754.806944444445, 23754.808333333334, 23754.80972222222, 23754.81111111111, 23754.8125, 23754.81388888889, 23754.81527777778, 23754.816666666666, 23754.818055555555, 23754.819444444445, 23754.820833333335, 23754.82222222222, 23754.82361111111, 23754.825, 23754.82638888889, 23754.827777777777, 23754.829166666666, 23754.830555555556, 23754.831944444446, 23754.833333333332, 23754.834722222222, 23754.83611111111, 23754.8375, 23754.838888888888, 23754.840277777777, 23754.841666666667, 23754.843055555557, 23754.844444444443, 23754.845833333333, 23754.847222222223, 23754.848611111112, 23754.85, 23754.85138888889, 23754.852777777778, 23754.854166666668, 23754.855555555554, 23754.856944444444, 23754.858333333334, 23754.859722222223, 23754.86111111111, 23754.8625, 23754.86388888889, 23754.86527777778, 23754.866666666665, 23754.868055555555, 23754.869444444445, 23754.870833333334, 23754.87222222222, 23754.87361111111, 23754.875, 23754.87638888889, 23754.87777777778, 23754.879166666666, 23754.880555555555, 23754.881944444445, 23754.883333333335, 23754.88472222222, 23754.88611111111, 23754.8875, 23754.88888888889, 23754.890277777777, 23754.891666666666, 23754.893055555556, 23754.894444444446, 23754.895833333332, 23754.897222222222, 23754.89861111111, 23754.9, 23754.901388888888, 23754.902777777777, 23754.904166666667, 23754.905555555557, 23754.906944444443, 23754.908333333333, 23754.909722222223, 23754.911111111112, 23754.9125, 23754.91388888889, 23754.915277777778, 23754.916666666668, 23754.918055555554, 23754.919444444444, 23754.920833333334, 23754.922222222223, 23754.92361111111, 23754.925, 23754.92638888889, 23754.92777777778, 23754.929166666665, 23754.930555555555, 23754.931944444445, 23754.933333333334, 23754.93472222222, 23754.93611111111, 23754.9375, 23754.93888888889, 23754.94027777778, 23754.941666666666, 23754.943055555555, 23754.944444444445, 23754.945833333335, 23754.94722222222, 23754.94861111111, 23754.95, 23754.95138888889, 23754.952777777777, 23754.954166666666, 23754.955555555556, 23754.956944444446, 23754.958333333332, 23754.959722222222, 23754.96111111111, 23754.9625, 23754.963888888888, 23754.965277777777, 23754.966666666667, 23754.968055555557, 23754.969444444443, 23754.970833333333, 23754.972222222223, 23754.973611111112, 23754.975, 23754.97638888889, 23754.977777777778, 23754.979166666668, 23754.980555555554, 23754.981944444444, 23754.983333333334, 23754.984722222223, 23754.98611111111, 23754.9875, 23754.98888888889, 23754.99027777778, 23754.991666666665, 23754.993055555555, 23754.994444444445, 23754.995833333334, 23754.99722222222, 23754.99861111111, 23755.0, 23755.00138888889, 23755.00277777778, 23755.004166666666, 23755.005555555555, 23755.006944444445, 23755.008333333335, 23755.00972222222, 23755.01111111111, 23755.0125, 23755.01388888889, 23755.015277777777, 23755.016666666666, 23755.018055555556, 23755.019444444446, 23755.020833333332, 23755.022222222222, 23755.02361111111, 23755.025, 23755.026388888888, 23755.027777777777, 23755.029166666667, 23755.030555555557, 23755.031944444443, 23755.033333333333, 23755.034722222223, 23755.036111111112, 23755.0375, 23755.03888888889, 23755.040277777778, 23755.041666666668, 23755.043055555554, 23755.044444444444, 23755.045833333334, 23755.047222222223, 23755.04861111111, 23755.05, 23755.05138888889, 23755.05277777778, 23755.054166666665, 23755.055555555555, 23755.056944444445, 23755.058333333334, 23755.05972222222, 23755.06111111111, 23755.0625, 23755.06388888889, 23755.06527777778, 23755.066666666666, 23755.068055555555, 23755.069444444445, 23755.070833333335, 23755.07222222222, 23755.07361111111, 23755.075, 23755.07638888889, 23755.077777777777, 23755.079166666666, 23755.080555555556, 23755.081944444446, 23755.083333333332, 23755.084722222222, 23755.08611111111, 23755.0875, 23755.088888888888, 23755.090277777777, 23755.091666666667, 23755.093055555557, 23755.094444444443, 23755.095833333333, 23755.097222222223, 23755.098611111112, 23755.1, 23755.10138888889, 23755.102777777778, 23755.104166666668, 23755.105555555554, 23755.106944444444, 23755.108333333334, 23755.109722222223, 23755.11111111111, 23755.1125, 23755.11388888889, 23755.11527777778, 23755.116666666665, 23755.118055555555, 23755.119444444445, 23755.120833333334, 23755.12222222222, 23755.12361111111, 23755.125, 23755.12638888889, 23755.12777777778, 23755.129166666666, 23755.130555555555, 23755.131944444445, 23755.133333333335, 23755.13472222222, 23755.13611111111, 23755.1375, 23755.13888888889, 23755.140277777777, 23755.141666666666, 23755.143055555556, 23755.144444444446, 23755.145833333332, 23755.147222222222, 23755.14861111111, 23755.15, 23755.151388888888, 23755.152777777777, 23755.154166666667, 23755.155555555557, 23755.156944444443, 23755.158333333333, 23755.159722222223, 23755.161111111112, 23755.1625, 23755.16388888889, 23755.165277777778, 23755.166666666668, 23755.168055555554, 23755.169444444444, 23755.170833333334, 23755.172222222223, 23755.17361111111, 23755.175, 23755.17638888889, 23755.17777777778, 23755.179166666665, 23755.180555555555, 23755.181944444445, 23755.183333333334, 23755.18472222222, 23755.18611111111, 23755.1875, 23755.18888888889, 23755.19027777778, 23755.191666666666, 23755.193055555555, 23755.194444444445, 23755.195833333335, 23755.19722222222, 23755.19861111111, 23755.2, 23755.20138888889, 23755.202777777777, 23755.204166666666, 23755.205555555556, 23755.206944444446, 23755.208333333332, 23755.209722222222, 23755.21111111111, 23755.2125, 23755.213888888888, 23755.215277777777, 23755.216666666667, 23755.218055555557, 23755.219444444443, 23755.220833333333, 23755.222222222223, 23755.223611111112, 23755.225, 23755.22638888889, 23755.227777777778, 23755.229166666668, 23755.230555555554, 23755.231944444444, 23755.233333333334, 23755.234722222223, 23755.23611111111, 23755.2375, 23755.23888888889, 23755.24027777778, 23755.241666666665, 23755.243055555555, 23755.244444444445, 23755.245833333334, 23755.24722222222, 23755.24861111111, 23755.25, 23755.25138888889, 23755.25277777778, 23755.254166666666, 23755.255555555555, 23755.256944444445, 23755.258333333335, 23755.25972222222, 23755.26111111111, 23755.2625, 23755.26388888889, 23755.265277777777, 23755.266666666666, 23755.268055555556, 23755.269444444446, 23755.270833333332, 23755.272222222222, 23755.27361111111, 23755.275, 23755.276388888888, 23755.277777777777, 23755.279166666667, 23755.280555555557, 23755.281944444443, 23755.283333333333, 23755.284722222223, 23755.286111111112, 23755.2875, 23755.28888888889, 23755.290277777778, 23755.291666666668, 23755.293055555554, 23755.294444444444, 23755.295833333334, 23755.297222222223, 23755.29861111111, 23755.3, 23755.30138888889, 23755.30277777778, 23755.304166666665, 23755.305555555555, 23755.306944444445, 23755.308333333334, 23755.30972222222, 23755.31111111111, 23755.3125, 23755.31388888889, 23755.31527777778, 23755.316666666666, 23755.318055555555, 23755.319444444445, 23755.320833333335, 23755.32222222222, 23755.32361111111, 23755.325, 23755.32638888889, 23755.327777777777, 23755.329166666666, 23755.330555555556, 23755.331944444446, 23755.333333333332, 23755.334722222222, 23755.33611111111, 23755.3375, 23755.338888888888, 23755.340277777777, 23755.341666666667, 23755.343055555557, 23755.344444444443, 23755.345833333333, 23755.347222222223, 23755.348611111112, 23755.35, 23755.35138888889, 23755.352777777778, 23755.354166666668, 23755.355555555554, 23755.356944444444, 23755.358333333334, 23755.359722222223, 23755.36111111111, 23755.3625, 23755.36388888889, 23755.36527777778, 23755.366666666665, 23755.368055555555, 23755.369444444445, 23755.370833333334, 23755.37222222222, 23755.37361111111, 23755.375, 23755.37638888889, 23755.37777777778, 23755.379166666666, 23755.380555555555, 23755.381944444445, 23755.383333333335, 23755.38472222222, 23755.38611111111, 23755.3875, 23755.38888888889, 23755.390277777777, 23755.391666666666, 23755.393055555556, 23755.394444444446, 23755.395833333332, 23755.397222222222, 23755.39861111111, 23755.4, 23755.401388888888, 23755.402777777777, 23755.404166666667, 23755.405555555557, 23755.406944444443, 23755.408333333333, 23755.409722222223, 23755.411111111112, 23755.4125, 23755.41388888889, 23755.415277777778, 23755.416666666668, 23755.418055555554, 23755.419444444444, 23755.420833333334, 23755.422222222223, 23755.42361111111, 23755.425, 23755.42638888889, 23755.42777777778, 23755.429166666665, 23755.430555555555, 23755.431944444445, 23755.433333333334, 23755.43472222222, 23755.43611111111, 23755.4375, 23755.43888888889, 23755.44027777778, 23755.441666666666, 23755.443055555555, 23755.444444444445, 23755.445833333335, 23755.44722222222, 23755.44861111111, 23755.45, 23755.45138888889, 23755.452777777777, 23755.454166666666, 23755.455555555556, 23755.456944444446, 23755.458333333332, 23755.459722222222, 23755.46111111111, 23755.4625, 23755.463888888888, 23755.465277777777, 23755.466666666667, 23755.468055555557, 23755.469444444443, 23755.470833333333, 23755.472222222223, 23755.473611111112, 23755.475, 23755.47638888889, 23755.477777777778, 23755.479166666668, 23755.480555555554, 23755.481944444444, 23755.483333333334, 23755.484722222223, 23755.48611111111, 23755.4875, 23755.48888888889, 23755.49027777778, 23755.491666666665, 23755.493055555555, 23755.494444444445, 23755.495833333334, 23755.49722222222, 23755.49861111111, 23755.5, 23755.50138888889, 23755.50277777778, 23755.504166666666, 23755.505555555555, 23755.506944444445, 23755.508333333335, 23755.50972222222, 23755.51111111111, 23755.5125, 23755.51388888889, 23755.515277777777, 23755.516666666666, 23755.518055555556, 23755.519444444446, 23755.520833333332, 23755.522222222222, 23755.52361111111, 23755.525, 23755.526388888888, 23755.527777777777, 23755.529166666667, 23755.530555555557, 23755.531944444443, 23755.533333333333, 23755.534722222223, 23755.536111111112, 23755.5375, 23755.53888888889, 23755.540277777778, 23755.541666666668, 23755.543055555554, 23755.544444444444, 23755.545833333334, 23755.547222222223, 23755.54861111111, 23755.55, 23755.55138888889, 23755.55277777778, 23755.554166666665, 23755.555555555555, 23755.556944444445, 23755.558333333334, 23755.55972222222, 23755.56111111111, 23755.5625, 23755.56388888889, 23755.56527777778, 23755.566666666666, 23755.568055555555, 23755.569444444445, 23755.570833333335, 23755.57222222222, 23755.57361111111, 23755.575, 23755.57638888889, 23755.577777777777, 23755.579166666666, 23755.580555555556, 23755.581944444446, 23755.583333333332, 23755.584722222222, 23755.58611111111, 23755.5875, 23755.588888888888, 23755.590277777777, 23755.591666666667, 23755.593055555557, 23755.594444444443, 23755.595833333333, 23755.597222222223, 23755.598611111112, 23755.6, 23755.60138888889, 23755.602777777778, 23755.604166666668, 23755.605555555554, 23755.606944444444, 23755.608333333334, 23755.609722222223, 23755.61111111111, 23755.6125, 23755.61388888889, 23755.61527777778, 23755.616666666665, 23755.618055555555, 23755.619444444445, 23755.620833333334, 23755.62222222222, 23755.62361111111, 23755.625, 23755.62638888889, 23755.62777777778, 23755.629166666666, 23755.630555555555, 23755.631944444445, 23755.633333333335, 23755.63472222222, 23755.63611111111, 23755.6375, 23755.63888888889, 23755.640277777777, 23755.641666666666, 23755.643055555556, 23755.644444444446, 23755.645833333332, 23755.647222222222, 23755.64861111111, 23755.65, 23755.651388888888, 23755.652777777777, 23755.654166666667, 23755.655555555557, 23755.656944444443, 23755.658333333333, 23755.659722222223, 23755.661111111112, 23755.6625, 23755.66388888889, 23755.665277777778, 23755.666666666668, 23755.668055555554, 23755.669444444444, 23755.670833333334, 23755.672222222223, 23755.67361111111, 23755.675, 23755.67638888889, 23755.67777777778, 23755.679166666665, 23755.680555555555, 23755.681944444445, 23755.683333333334, 23755.68472222222, 23755.68611111111, 23755.6875, 23755.68888888889, 23755.69027777778, 23755.691666666666, 23755.693055555555, 23755.694444444445, 23755.695833333335, 23755.69722222222, 23755.69861111111, 23755.7, 23755.70138888889, 23755.702777777777, 23755.704166666666, 23755.705555555556, 23755.706944444446, 23755.708333333332, 23755.709722222222, 23755.71111111111, 23755.7125, 23755.713888888888, 23755.715277777777, 23755.716666666667, 23755.718055555557, 23755.719444444443, 23755.720833333333, 23755.722222222223, 23755.723611111112, 23755.725, 23755.72638888889, 23755.727777777778, 23755.729166666668, 23755.730555555554, 23755.731944444444, 23755.733333333334, 23755.734722222223, 23755.73611111111, 23755.7375, 23755.73888888889, 23755.74027777778, 23755.741666666665, 23755.743055555555, 23755.744444444445, 23755.745833333334, 23755.74722222222, 23755.74861111111, 23755.75, 23755.75138888889, 23755.75277777778, 23755.754166666666, 23755.755555555555, 23755.756944444445, 23755.758333333335, 23755.75972222222, 23755.76111111111, 23755.7625, 23755.76388888889, 23755.765277777777, 23755.766666666666, 23755.768055555556, 23755.769444444446, 23755.770833333332, 23755.772222222222, 23755.77361111111, 23755.775, 23755.776388888888, 23755.777777777777, 23755.779166666667, 23755.780555555557, 23755.781944444443, 23755.783333333333, 23755.784722222223, 23755.786111111112, 23755.7875, 23755.78888888889, 23755.790277777778, 23755.791666666668, 23755.793055555554, 23755.794444444444, 23755.795833333334, 23755.797222222223, 23755.79861111111, 23755.8, 23755.80138888889, 23755.80277777778, 23755.804166666665, 23755.805555555555, 23755.806944444445, 23755.808333333334, 23755.80972222222, 23755.81111111111, 23755.8125, 23755.81388888889, 23755.81527777778, 23755.816666666666, 23755.818055555555, 23755.819444444445, 23755.820833333335, 23755.82222222222, 23755.82361111111, 23755.825, 23755.82638888889, 23755.827777777777, 23755.829166666666, 23755.830555555556, 23755.831944444446, 23755.833333333332, 23755.834722222222, 23755.83611111111, 23755.8375, 23755.838888888888, 23755.840277777777, 23755.841666666667, 23755.843055555557, 23755.844444444443, 23755.845833333333, 23755.847222222223, 23755.848611111112, 23755.85, 23755.85138888889, 23755.852777777778, 23755.854166666668, 23755.855555555554, 23755.856944444444, 23755.858333333334, 23755.859722222223, 23755.86111111111, 23755.8625, 23755.86388888889, 23755.86527777778, 23755.866666666665, 23755.868055555555, 23755.869444444445, 23755.870833333334, 23755.87222222222, 23755.87361111111, 23755.875, 23755.87638888889, 23755.87777777778, 23755.879166666666, 23755.880555555555, 23755.881944444445, 23755.883333333335, 23755.88472222222, 23755.88611111111, 23755.8875, 23755.88888888889, 23755.890277777777, 23755.891666666666, 23755.893055555556, 23755.894444444446, 23755.895833333332, 23755.897222222222, 23755.89861111111, 23755.9, 23755.901388888888, 23755.902777777777, 23755.904166666667, 23755.905555555557, 23755.906944444443, 23755.908333333333, 23755.909722222223, 23755.911111111112, 23755.9125, 23755.91388888889, 23755.915277777778, 23755.916666666668, 23755.918055555554, 23755.919444444444, 23755.920833333334, 23755.922222222223, 23755.92361111111, 23755.925, 23755.92638888889, 23755.92777777778, 23755.929166666665, 23755.930555555555, 23755.931944444445, 23755.933333333334, 23755.93472222222, 23755.93611111111, 23755.9375, 23755.93888888889, 23755.94027777778, 23755.941666666666, 23755.943055555555, 23755.944444444445, 23755.945833333335, 23755.94722222222, 23755.94861111111, 23755.95, 23755.95138888889, 23755.952777777777, 23755.954166666666, 23755.955555555556, 23755.956944444446, 23755.958333333332, 23755.959722222222, 23755.96111111111, 23755.9625, 23755.963888888888, 23755.965277777777, 23755.966666666667, 23755.968055555557, 23755.969444444443, 23755.970833333333, 23755.972222222223, 23755.973611111112, 23755.975, 23755.97638888889, 23755.977777777778, 23755.979166666668, 23755.980555555554, 23755.981944444444, 23755.983333333334, 23755.984722222223, 23755.98611111111, 23755.9875, 23755.98888888889, 23755.99027777778, 23755.991666666665, 23755.993055555555, 23755.994444444445, 23755.995833333334, 23755.99722222222, 23755.99861111111, 23756.0, 23756.00138888889, 23756.00277777778, 23756.004166666666, 23756.005555555555, 23756.006944444445, 23756.008333333335, 23756.00972222222, 23756.01111111111, 23756.0125, 23756.01388888889, 23756.015277777777, 23756.016666666666, 23756.018055555556, 23756.019444444446, 23756.020833333332, 23756.022222222222, 23756.02361111111, 23756.025, 23756.026388888888, 23756.027777777777, 23756.029166666667, 23756.030555555557, 23756.031944444443, 23756.033333333333, 23756.034722222223, 23756.036111111112, 23756.0375, 23756.03888888889, 23756.040277777778, 23756.041666666668, 23756.043055555554, 23756.044444444444, 23756.045833333334, 23756.047222222223, 23756.04861111111, 23756.05, 23756.05138888889, 23756.05277777778, 23756.054166666665, 23756.055555555555, 23756.056944444445, 23756.058333333334, 23756.05972222222, 23756.06111111111, 23756.0625, 23756.06388888889, 23756.06527777778, 23756.066666666666, 23756.068055555555, 23756.069444444445, 23756.070833333335, 23756.07222222222, 23756.07361111111, 23756.075, 23756.07638888889, 23756.077777777777, 23756.079166666666, 23756.080555555556, 23756.081944444446, 23756.083333333332, 23756.084722222222, 23756.08611111111, 23756.0875, 23756.088888888888, 23756.090277777777, 23756.091666666667, 23756.093055555557, 23756.094444444443, 23756.095833333333, 23756.097222222223, 23756.098611111112, 23756.1, 23756.10138888889, 23756.102777777778, 23756.104166666668, 23756.105555555554, 23756.106944444444, 23756.108333333334, 23756.109722222223, 23756.11111111111, 23756.1125, 23756.11388888889, 23756.11527777778, 23756.116666666665, 23756.118055555555, 23756.119444444445, 23756.120833333334, 23756.12222222222, 23756.12361111111, 23756.125, 23756.12638888889, 23756.12777777778, 23756.129166666666, 23756.130555555555, 23756.131944444445, 23756.133333333335, 23756.13472222222, 23756.13611111111, 23756.1375, 23756.13888888889, 23756.140277777777, 23756.141666666666, 23756.143055555556, 23756.144444444446, 23756.145833333332, 23756.147222222222, 23756.14861111111, 23756.15, 23756.151388888888, 23756.152777777777, 23756.154166666667, 23756.155555555557, 23756.156944444443, 23756.158333333333, 23756.159722222223, 23756.161111111112, 23756.1625, 23756.16388888889, 23756.165277777778, 23756.166666666668, 23756.168055555554, 23756.169444444444, 23756.170833333334, 23756.172222222223, 23756.17361111111, 23756.175, 23756.17638888889, 23756.17777777778, 23756.179166666665, 23756.180555555555, 23756.181944444445, 23756.183333333334, 23756.18472222222, 23756.18611111111, 23756.1875, 23756.18888888889, 23756.19027777778, 23756.191666666666, 23756.193055555555, 23756.194444444445, 23756.195833333335, 23756.19722222222, 23756.19861111111, 23756.2, 23756.20138888889, 23756.202777777777, 23756.204166666666, 23756.205555555556, 23756.206944444446, 23756.208333333332, 23756.209722222222, 23756.21111111111, 23756.2125, 23756.213888888888, 23756.215277777777, 23756.216666666667, 23756.218055555557, 23756.219444444443, 23756.220833333333, 23756.222222222223, 23756.223611111112, 23756.225, 23756.22638888889, 23756.227777777778, 23756.229166666668, 23756.230555555554, 23756.231944444444, 23756.233333333334, 23756.234722222223, 23756.23611111111, 23756.2375, 23756.23888888889, 23756.24027777778, 23756.241666666665, 23756.243055555555, 23756.244444444445, 23756.245833333334, 23756.24722222222, 23756.24861111111, 23756.25, 23756.25138888889, 23756.25277777778, 23756.254166666666, 23756.255555555555, 23756.256944444445, 23756.258333333335, 23756.25972222222, 23756.26111111111, 23756.2625, 23756.26388888889, 23756.265277777777, 23756.266666666666, 23756.268055555556, 23756.269444444446, 23756.270833333332, 23756.272222222222, 23756.27361111111, 23756.275, 23756.276388888888, 23756.277777777777, 23756.279166666667, 23756.280555555557, 23756.281944444443, 23756.283333333333, 23756.284722222223, 23756.286111111112, 23756.2875, 23756.28888888889, 23756.290277777778, 23756.291666666668, 23756.293055555554, 23756.294444444444, 23756.295833333334, 23756.297222222223, 23756.29861111111, 23756.3, 23756.30138888889, 23756.30277777778, 23756.304166666665, 23756.305555555555, 23756.306944444445, 23756.308333333334, 23756.30972222222, 23756.31111111111, 23756.3125, 23756.31388888889, 23756.31527777778, 23756.316666666666, 23756.318055555555, 23756.319444444445, 23756.320833333335, 23756.32222222222, 23756.32361111111, 23756.325, 23756.32638888889, 23756.327777777777, 23756.329166666666, 23756.330555555556, 23756.331944444446, 23756.333333333332, 23756.334722222222, 23756.33611111111, 23756.3375, 23756.338888888888, 23756.340277777777, 23756.341666666667, 23756.343055555557, 23756.344444444443, 23756.345833333333, 23756.347222222223, 23756.348611111112, 23756.35, 23756.35138888889, 23756.352777777778, 23756.354166666668, 23756.355555555554, 23756.356944444444, 23756.358333333334, 23756.359722222223, 23756.36111111111, 23756.3625, 23756.36388888889, 23756.36527777778, 23756.366666666665, 23756.368055555555, 23756.369444444445, 23756.370833333334, 23756.37222222222, 23756.37361111111, 23756.375, 23756.37638888889, 23756.37777777778, 23756.379166666666, 23756.380555555555, 23756.381944444445, 23756.383333333335, 23756.38472222222, 23756.38611111111, 23756.3875, 23756.38888888889, 23756.390277777777, 23756.391666666666, 23756.393055555556, 23756.394444444446, 23756.395833333332, 23756.397222222222, 23756.39861111111, 23756.4, 23756.401388888888, 23756.402777777777, 23756.404166666667, 23756.405555555557, 23756.406944444443, 23756.408333333333, 23756.409722222223, 23756.411111111112, 23756.4125, 23756.41388888889, 23756.415277777778, 23756.416666666668, 23756.418055555554, 23756.419444444444, 23756.420833333334, 23756.422222222223, 23756.42361111111, 23756.425, 23756.42638888889, 23756.42777777778, 23756.429166666665, 23756.430555555555, 23756.431944444445, 23756.433333333334, 23756.43472222222, 23756.43611111111, 23756.4375, 23756.43888888889, 23756.44027777778, 23756.441666666666, 23756.443055555555, 23756.444444444445, 23756.445833333335, 23756.44722222222, 23756.44861111111, 23756.45, 23756.45138888889, 23756.452777777777, 23756.454166666666, 23756.455555555556, 23756.456944444446, 23756.458333333332, 23756.459722222222, 23756.46111111111, 23756.4625, 23756.463888888888, 23756.465277777777, 23756.466666666667, 23756.468055555557, 23756.469444444443, 23756.470833333333, 23756.472222222223, 23756.473611111112, 23756.475, 23756.47638888889, 23756.477777777778, 23756.479166666668, 23756.480555555554, 23756.481944444444, 23756.483333333334, 23756.484722222223, 23756.48611111111, 23756.4875, 23756.48888888889, 23756.49027777778, 23756.491666666665, 23756.493055555555, 23756.494444444445, 23756.495833333334, 23756.49722222222, 23756.49861111111, 23756.5, 23756.50138888889, 23756.50277777778, 23756.504166666666, 23756.505555555555, 23756.506944444445, 23756.508333333335, 23756.50972222222, 23756.51111111111, 23756.5125, 23756.51388888889, 23756.515277777777, 23756.516666666666, 23756.518055555556, 23756.519444444446, 23756.520833333332, 23756.522222222222, 23756.52361111111, 23756.525, 23756.526388888888, 23756.527777777777, 23756.529166666667, 23756.530555555557, 23756.531944444443, 23756.533333333333, 23756.534722222223, 23756.536111111112, 23756.5375, 23756.53888888889, 23756.540277777778, 23756.541666666668, 23756.543055555554, 23756.544444444444, 23756.545833333334, 23756.547222222223, 23756.54861111111, 23756.55, 23756.55138888889, 23756.55277777778, 23756.554166666665, 23756.555555555555, 23756.556944444445, 23756.558333333334, 23756.55972222222, 23756.56111111111, 23756.5625, 23756.56388888889, 23756.56527777778, 23756.566666666666, 23756.568055555555, 23756.569444444445, 23756.570833333335, 23756.57222222222, 23756.57361111111, 23756.575, 23756.57638888889, 23756.577777777777, 23756.579166666666, 23756.580555555556, 23756.581944444446, 23756.583333333332, 23756.584722222222, 23756.58611111111, 23756.5875, 23756.588888888888, 23756.590277777777, 23756.591666666667, 23756.593055555557, 23756.594444444443, 23756.595833333333, 23756.597222222223, 23756.598611111112, 23756.6, 23756.60138888889, 23756.602777777778, 23756.604166666668, 23756.605555555554, 23756.606944444444, 23756.608333333334, 23756.609722222223, 23756.61111111111, 23756.6125, 23756.61388888889, 23756.61527777778, 23756.616666666665, 23756.618055555555, 23756.619444444445, 23756.620833333334, 23756.62222222222, 23756.62361111111, 23756.625, 23756.62638888889, 23756.62777777778, 23756.629166666666, 23756.630555555555, 23756.631944444445, 23756.633333333335, 23756.63472222222, 23756.63611111111, 23756.6375, 23756.63888888889, 23756.640277777777, 23756.641666666666, 23756.643055555556, 23756.644444444446, 23756.645833333332, 23756.647222222222, 23756.64861111111, 23756.65, 23756.651388888888, 23756.652777777777, 23756.654166666667, 23756.655555555557, 23756.656944444443, 23756.658333333333, 23756.659722222223, 23756.661111111112, 23756.6625, 23756.66388888889, 23756.665277777778, 23756.666666666668, 23756.668055555554, 23756.669444444444, 23756.670833333334, 23756.672222222223, 23756.67361111111, 23756.675, 23756.67638888889, 23756.67777777778, 23756.679166666665, 23756.680555555555, 23756.681944444445, 23756.683333333334, 23756.68472222222, 23756.68611111111, 23756.6875, 23756.68888888889, 23756.69027777778, 23756.691666666666, 23756.693055555555, 23756.694444444445, 23756.695833333335, 23756.69722222222, 23756.69861111111, 23756.7, 23756.70138888889, 23756.702777777777, 23756.704166666666, 23756.705555555556, 23756.706944444446, 23756.708333333332, 23756.709722222222, 23756.71111111111, 23756.7125, 23756.713888888888, 23756.715277777777, 23756.716666666667, 23756.718055555557, 23756.719444444443, 23756.720833333333, 23756.722222222223, 23756.723611111112, 23756.725, 23756.72638888889, 23756.727777777778, 23756.729166666668, 23756.730555555554, 23756.731944444444, 23756.733333333334, 23756.734722222223, 23756.73611111111, 23756.7375, 23756.73888888889, 23756.74027777778, 23756.741666666665, 23756.743055555555, 23756.744444444445, 23756.745833333334, 23756.74722222222, 23756.74861111111, 23756.75, 23756.75138888889, 23756.75277777778, 23756.754166666666, 23756.755555555555, 23756.756944444445, 23756.758333333335, 23756.75972222222, 23756.76111111111, 23756.7625, 23756.76388888889, 23756.765277777777, 23756.766666666666, 23756.768055555556, 23756.769444444446, 23756.770833333332, 23756.772222222222, 23756.77361111111, 23756.775, 23756.776388888888, 23756.777777777777, 23756.779166666667, 23756.780555555557, 23756.781944444443, 23756.783333333333, 23756.784722222223, 23756.786111111112, 23756.7875, 23756.78888888889, 23756.790277777778, 23756.791666666668, 23756.793055555554, 23756.794444444444, 23756.795833333334, 23756.797222222223, 23756.79861111111, 23756.8, 23756.80138888889, 23756.80277777778, 23756.804166666665, 23756.805555555555, 23756.806944444445, 23756.808333333334, 23756.80972222222, 23756.81111111111, 23756.8125, 23756.81388888889, 23756.81527777778, 23756.816666666666, 23756.818055555555, 23756.819444444445, 23756.820833333335, 23756.82222222222, 23756.82361111111, 23756.825, 23756.82638888889, 23756.827777777777, 23756.829166666666, 23756.830555555556, 23756.831944444446, 23756.833333333332, 23756.834722222222, 23756.83611111111, 23756.8375, 23756.838888888888, 23756.840277777777, 23756.841666666667, 23756.843055555557, 23756.844444444443, 23756.845833333333, 23756.847222222223, 23756.848611111112, 23756.85, 23756.85138888889, 23756.852777777778, 23756.854166666668, 23756.855555555554, 23756.856944444444, 23756.858333333334, 23756.859722222223, 23756.86111111111, 23756.8625, 23756.86388888889, 23756.86527777778, 23756.866666666665, 23756.868055555555, 23756.869444444445, 23756.870833333334, 23756.87222222222, 23756.87361111111, 23756.875, 23756.87638888889, 23756.87777777778, 23756.879166666666, 23756.880555555555, 23756.881944444445, 23756.883333333335, 23756.88472222222, 23756.88611111111, 23756.8875, 23756.88888888889, 23756.890277777777, 23756.891666666666, 23756.893055555556, 23756.894444444446, 23756.895833333332, 23756.897222222222, 23756.89861111111, 23756.9, 23756.901388888888, 23756.902777777777, 23756.904166666667, 23756.905555555557, 23756.906944444443, 23756.908333333333, 23756.909722222223, 23756.911111111112, 23756.9125, 23756.91388888889, 23756.915277777778, 23756.916666666668, 23756.918055555554, 23756.919444444444, 23756.920833333334, 23756.922222222223, 23756.92361111111, 23756.925, 23756.92638888889, 23756.92777777778, 23756.929166666665, 23756.930555555555, 23756.931944444445, 23756.933333333334, 23756.93472222222, 23756.93611111111, 23756.9375, 23756.93888888889, 23756.94027777778, 23756.941666666666, 23756.943055555555, 23756.944444444445, 23756.945833333335, 23756.94722222222, 23756.94861111111, 23756.95, 23756.95138888889, 23756.952777777777, 23756.954166666666, 23756.955555555556, 23756.956944444446, 23756.958333333332, 23756.959722222222, 23756.96111111111, 23756.9625, 23756.963888888888, 23756.965277777777, 23756.966666666667, 23756.968055555557, 23756.969444444443, 23756.970833333333, 23756.972222222223, 23756.973611111112, 23756.975, 23756.97638888889, 23756.977777777778, 23756.979166666668, 23756.980555555554, 23756.981944444444, 23756.983333333334, 23756.984722222223, 23756.98611111111, 23756.9875, 23756.98888888889, 23756.99027777778, 23756.991666666665, 23756.993055555555, 23756.994444444445, 23756.995833333334, 23756.99722222222, 23756.99861111111, 23757.0, 23757.00138888889, 23757.00277777778, 23757.004166666666, 23757.005555555555, 23757.006944444445, 23757.008333333335, 23757.00972222222, 23757.01111111111, 23757.0125, 23757.01388888889, 23757.015277777777, 23757.016666666666, 23757.018055555556, 23757.019444444446, 23757.020833333332, 23757.022222222222, 23757.02361111111, 23757.025, 23757.026388888888, 23757.027777777777, 23757.029166666667, 23757.030555555557, 23757.031944444443, 23757.033333333333, 23757.034722222223, 23757.036111111112, 23757.0375, 23757.03888888889, 23757.040277777778, 23757.041666666668, 23757.043055555554, 23757.044444444444, 23757.045833333334, 23757.047222222223, 23757.04861111111, 23757.05, 23757.05138888889, 23757.05277777778, 23757.054166666665, 23757.055555555555, 23757.056944444445, 23757.058333333334, 23757.05972222222, 23757.06111111111, 23757.0625, 23757.06388888889, 23757.06527777778, 23757.066666666666, 23757.068055555555, 23757.069444444445, 23757.070833333335, 23757.07222222222, 23757.07361111111, 23757.075, 23757.07638888889, 23757.077777777777, 23757.079166666666, 23757.080555555556, 23757.081944444446, 23757.083333333332, 23757.084722222222, 23757.08611111111, 23757.0875, 23757.088888888888, 23757.090277777777, 23757.091666666667, 23757.093055555557, 23757.094444444443, 23757.095833333333, 23757.097222222223, 23757.098611111112, 23757.1, 23757.10138888889, 23757.102777777778, 23757.104166666668, 23757.105555555554, 23757.106944444444, 23757.108333333334, 23757.109722222223, 23757.11111111111, 23757.1125, 23757.11388888889, 23757.11527777778, 23757.116666666665, 23757.118055555555, 23757.119444444445, 23757.120833333334, 23757.12222222222, 23757.12361111111, 23757.125, 23757.12638888889, 23757.12777777778, 23757.129166666666, 23757.130555555555, 23757.131944444445, 23757.133333333335, 23757.13472222222, 23757.13611111111, 23757.1375, 23757.13888888889, 23757.140277777777, 23757.141666666666, 23757.143055555556, 23757.144444444446, 23757.145833333332, 23757.147222222222, 23757.14861111111, 23757.15, 23757.151388888888, 23757.152777777777, 23757.154166666667, 23757.155555555557, 23757.156944444443, 23757.158333333333, 23757.159722222223, 23757.161111111112, 23757.1625, 23757.16388888889, 23757.165277777778, 23757.166666666668, 23757.168055555554, 23757.169444444444, 23757.170833333334, 23757.172222222223, 23757.17361111111, 23757.175, 23757.17638888889, 23757.17777777778, 23757.179166666665, 23757.180555555555, 23757.181944444445, 23757.183333333334, 23757.18472222222, 23757.18611111111, 23757.1875, 23757.18888888889, 23757.19027777778, 23757.191666666666, 23757.193055555555, 23757.194444444445, 23757.195833333335, 23757.19722222222, 23757.19861111111, 23757.2, 23757.20138888889, 23757.202777777777, 23757.204166666666, 23757.205555555556, 23757.206944444446, 23757.208333333332, 23757.209722222222, 23757.21111111111, 23757.2125, 23757.213888888888, 23757.215277777777, 23757.216666666667, 23757.218055555557, 23757.219444444443, 23757.220833333333, 23757.222222222223, 23757.223611111112, 23757.225, 23757.22638888889, 23757.227777777778, 23757.229166666668, 23757.230555555554, 23757.231944444444, 23757.233333333334, 23757.234722222223, 23757.23611111111, 23757.2375, 23757.23888888889, 23757.24027777778, 23757.241666666665, 23757.243055555555, 23757.244444444445, 23757.245833333334, 23757.24722222222, 23757.24861111111, 23757.25, 23757.25138888889, 23757.25277777778, 23757.254166666666, 23757.255555555555, 23757.256944444445, 23757.258333333335, 23757.25972222222, 23757.26111111111, 23757.2625, 23757.26388888889, 23757.265277777777, 23757.266666666666, 23757.268055555556, 23757.269444444446, 23757.270833333332, 23757.272222222222, 23757.27361111111, 23757.275, 23757.276388888888, 23757.277777777777, 23757.279166666667, 23757.280555555557, 23757.281944444443, 23757.283333333333, 23757.284722222223, 23757.286111111112, 23757.2875, 23757.28888888889, 23757.290277777778, 23757.291666666668, 23757.293055555554, 23757.294444444444, 23757.295833333334, 23757.297222222223, 23757.29861111111, 23757.3, 23757.30138888889, 23757.30277777778, 23757.304166666665, 23757.305555555555, 23757.306944444445, 23757.308333333334, 23757.30972222222, 23757.31111111111, 23757.3125, 23757.31388888889, 23757.31527777778, 23757.316666666666, 23757.318055555555, 23757.319444444445, 23757.320833333335, 23757.32222222222, 23757.32361111111, 23757.325, 23757.32638888889, 23757.327777777777, 23757.329166666666, 23757.330555555556, 23757.331944444446, 23757.333333333332, 23757.334722222222, 23757.33611111111, 23757.3375, 23757.338888888888, 23757.340277777777, 23757.341666666667, 23757.343055555557, 23757.344444444443, 23757.345833333333, 23757.347222222223, 23757.348611111112, 23757.35, 23757.35138888889, 23757.352777777778, 23757.354166666668, 23757.355555555554, 23757.356944444444, 23757.358333333334, 23757.359722222223, 23757.36111111111, 23757.3625, 23757.36388888889, 23757.36527777778, 23757.366666666665, 23757.368055555555, 23757.369444444445, 23757.370833333334, 23757.37222222222, 23757.37361111111, 23757.375, 23757.37638888889, 23757.37777777778, 23757.379166666666, 23757.380555555555, 23757.381944444445, 23757.383333333335, 23757.38472222222, 23757.38611111111, 23757.3875, 23757.38888888889, 23757.390277777777, 23757.391666666666, 23757.393055555556, 23757.394444444446, 23757.395833333332, 23757.397222222222, 23757.39861111111, 23757.4, 23757.401388888888, 23757.402777777777, 23757.404166666667, 23757.405555555557, 23757.406944444443, 23757.408333333333, 23757.409722222223, 23757.411111111112, 23757.4125, 23757.41388888889, 23757.415277777778, 23757.416666666668, 23757.418055555554, 23757.419444444444, 23757.420833333334, 23757.422222222223, 23757.42361111111, 23757.425, 23757.42638888889, 23757.42777777778, 23757.429166666665, 23757.430555555555, 23757.431944444445, 23757.433333333334, 23757.43472222222, 23757.43611111111, 23757.4375, 23757.43888888889, 23757.44027777778, 23757.441666666666, 23757.443055555555, 23757.444444444445, 23757.445833333335, 23757.44722222222, 23757.44861111111, 23757.45, 23757.45138888889, 23757.452777777777, 23757.454166666666, 23757.455555555556, 23757.456944444446, 23757.458333333332, 23757.459722222222, 23757.46111111111, 23757.4625, 23757.463888888888, 23757.465277777777, 23757.466666666667, 23757.468055555557, 23757.469444444443, 23757.470833333333, 23757.472222222223, 23757.473611111112, 23757.475, 23757.47638888889, 23757.477777777778, 23757.479166666668, 23757.480555555554, 23757.481944444444, 23757.483333333334, 23757.484722222223, 23757.48611111111, 23757.4875, 23757.48888888889, 23757.49027777778, 23757.491666666665, 23757.493055555555, 23757.494444444445, 23757.495833333334, 23757.49722222222, 23757.49861111111, 23757.5, 23757.50138888889, 23757.50277777778, 23757.504166666666, 23757.505555555555, 23757.506944444445, 23757.508333333335, 23757.50972222222, 23757.51111111111, 23757.5125, 23757.51388888889, 23757.515277777777, 23757.516666666666, 23757.518055555556, 23757.519444444446, 23757.520833333332, 23757.522222222222, 23757.52361111111, 23757.525, 23757.526388888888, 23757.527777777777, 23757.529166666667, 23757.530555555557, 23757.531944444443, 23757.533333333333, 23757.534722222223, 23757.536111111112, 23757.5375, 23757.53888888889, 23757.540277777778, 23757.541666666668, 23757.543055555554, 23757.544444444444, 23757.545833333334, 23757.547222222223, 23757.54861111111, 23757.55, 23757.55138888889, 23757.55277777778, 23757.554166666665, 23757.555555555555, 23757.556944444445, 23757.558333333334, 23757.55972222222, 23757.56111111111, 23757.5625, 23757.56388888889, 23757.56527777778, 23757.566666666666, 23757.568055555555, 23757.569444444445, 23757.570833333335, 23757.57222222222, 23757.57361111111, 23757.575, 23757.57638888889, 23757.577777777777, 23757.579166666666, 23757.580555555556, 23757.581944444446, 23757.583333333332, 23757.584722222222, 23757.58611111111, 23757.5875, 23757.588888888888, 23757.590277777777, 23757.591666666667, 23757.593055555557, 23757.594444444443, 23757.595833333333, 23757.597222222223, 23757.598611111112, 23757.6, 23757.60138888889, 23757.602777777778, 23757.604166666668, 23757.605555555554, 23757.606944444444, 23757.608333333334, 23757.609722222223, 23757.61111111111, 23757.6125, 23757.61388888889, 23757.61527777778, 23757.616666666665, 23757.618055555555, 23757.619444444445, 23757.620833333334, 23757.62222222222, 23757.62361111111, 23757.625, 23757.62638888889, 23757.62777777778, 23757.629166666666, 23757.630555555555, 23757.631944444445, 23757.633333333335, 23757.63472222222, 23757.63611111111, 23757.6375, 23757.63888888889, 23757.640277777777, 23757.641666666666, 23757.643055555556, 23757.644444444446, 23757.645833333332, 23757.647222222222, 23757.64861111111, 23757.65, 23757.651388888888, 23757.652777777777, 23757.654166666667, 23757.655555555557, 23757.656944444443, 23757.658333333333, 23757.659722222223, 23757.661111111112, 23757.6625, 23757.66388888889, 23757.665277777778, 23757.666666666668, 23757.668055555554, 23757.669444444444, 23757.670833333334, 23757.672222222223, 23757.67361111111, 23757.675, 23757.67638888889, 23757.67777777778, 23757.679166666665, 23757.680555555555, 23757.681944444445, 23757.683333333334, 23757.68472222222, 23757.68611111111, 23757.6875, 23757.68888888889, 23757.69027777778, 23757.691666666666, 23757.693055555555, 23757.694444444445, 23757.695833333335, 23757.69722222222, 23757.69861111111, 23757.7, 23757.70138888889, 23757.702777777777, 23757.704166666666, 23757.705555555556, 23757.706944444446, 23757.708333333332, 23757.709722222222, 23757.71111111111, 23757.7125, 23757.713888888888, 23757.715277777777, 23757.716666666667, 23757.718055555557, 23757.719444444443, 23757.720833333333, 23757.722222222223, 23757.723611111112, 23757.725, 23757.72638888889, 23757.727777777778, 23757.729166666668, 23757.730555555554, 23757.731944444444, 23757.733333333334, 23757.734722222223, 23757.73611111111, 23757.7375, 23757.73888888889, 23757.74027777778, 23757.741666666665, 23757.743055555555, 23757.744444444445, 23757.745833333334, 23757.74722222222, 23757.74861111111, 23757.75, 23757.75138888889, 23757.75277777778, 23757.754166666666, 23757.755555555555, 23757.756944444445, 23757.758333333335, 23757.75972222222, 23757.76111111111, 23757.7625, 23757.76388888889, 23757.765277777777, 23757.766666666666, 23757.768055555556, 23757.769444444446, 23757.770833333332, 23757.772222222222, 23757.77361111111, 23757.775, 23757.776388888888, 23757.777777777777, 23757.779166666667, 23757.780555555557, 23757.781944444443, 23757.783333333333, 23757.784722222223, 23757.786111111112, 23757.7875, 23757.78888888889, 23757.790277777778, 23757.791666666668, 23757.793055555554, 23757.794444444444, 23757.795833333334, 23757.797222222223, 23757.79861111111, 23757.8, 23757.80138888889, 23757.80277777778, 23757.804166666665, 23757.805555555555, 23757.806944444445, 23757.808333333334, 23757.80972222222, 23757.81111111111, 23757.8125, 23757.81388888889, 23757.81527777778, 23757.816666666666, 23757.818055555555, 23757.819444444445, 23757.820833333335, 23757.82222222222, 23757.82361111111, 23757.825, 23757.82638888889, 23757.827777777777, 23757.829166666666, 23757.830555555556, 23757.831944444446, 23757.833333333332, 23757.834722222222, 23757.83611111111, 23757.8375, 23757.838888888888, 23757.840277777777, 23757.841666666667, 23757.843055555557, 23757.844444444443, 23757.845833333333, 23757.847222222223, 23757.848611111112, 23757.85, 23757.85138888889, 23757.852777777778, 23757.854166666668, 23757.855555555554, 23757.856944444444, 23757.858333333334, 23757.859722222223, 23757.86111111111, 23757.8625, 23757.86388888889, 23757.86527777778, 23757.866666666665, 23757.868055555555, 23757.869444444445, 23757.870833333334, 23757.87222222222, 23757.87361111111, 23757.875, 23757.87638888889, 23757.87777777778, 23757.879166666666, 23757.880555555555, 23757.881944444445, 23757.883333333335, 23757.88472222222, 23757.88611111111, 23757.8875, 23757.88888888889, 23757.890277777777, 23757.891666666666, 23757.893055555556, 23757.894444444446, 23757.895833333332, 23757.897222222222, 23757.89861111111, 23757.9, 23757.901388888888, 23757.902777777777, 23757.904166666667, 23757.905555555557, 23757.906944444443, 23757.908333333333, 23757.909722222223, 23757.911111111112, 23757.9125, 23757.91388888889, 23757.915277777778, 23757.916666666668, 23757.918055555554, 23757.919444444444, 23757.920833333334, 23757.922222222223, 23757.92361111111, 23757.925, 23757.92638888889, 23757.92777777778, 23757.929166666665, 23757.930555555555, 23757.931944444445, 23757.933333333334, 23757.93472222222, 23757.93611111111, 23757.9375, 23757.93888888889, 23757.94027777778, 23757.941666666666, 23757.943055555555, 23757.944444444445, 23757.945833333335, 23757.94722222222, 23757.94861111111, 23757.95, 23757.95138888889, 23757.952777777777, 23757.954166666666, 23757.955555555556, 23757.956944444446, 23757.958333333332, 23757.959722222222, 23757.96111111111, 23757.9625, 23757.963888888888, 23757.965277777777, 23757.966666666667, 23757.968055555557, 23757.969444444443, 23757.970833333333, 23757.972222222223, 23757.973611111112, 23757.975, 23757.97638888889, 23757.977777777778, 23757.979166666668, 23757.980555555554, 23757.981944444444, 23757.983333333334, 23757.984722222223, 23757.98611111111, 23757.9875, 23757.98888888889, 23757.99027777778, 23757.991666666665, 23757.993055555555, 23757.994444444445, 23757.995833333334, 23757.99722222222, 23757.99861111111, 23758.0, 23758.00138888889, 23758.00277777778, 23758.004166666666, 23758.005555555555, 23758.006944444445, 23758.008333333335, 23758.00972222222, 23758.01111111111, 23758.0125, 23758.01388888889, 23758.015277777777, 23758.016666666666, 23758.018055555556, 23758.019444444446, 23758.020833333332, 23758.022222222222, 23758.02361111111, 23758.025, 23758.026388888888, 23758.027777777777, 23758.029166666667, 23758.030555555557, 23758.031944444443, 23758.033333333333, 23758.034722222223, 23758.036111111112, 23758.0375, 23758.03888888889, 23758.040277777778, 23758.041666666668, 23758.043055555554, 23758.044444444444, 23758.045833333334, 23758.047222222223, 23758.04861111111, 23758.05, 23758.05138888889, 23758.05277777778, 23758.054166666665, 23758.055555555555, 23758.056944444445, 23758.058333333334, 23758.05972222222, 23758.06111111111, 23758.0625, 23758.06388888889, 23758.06527777778, 23758.066666666666, 23758.068055555555, 23758.069444444445, 23758.070833333335, 23758.07222222222, 23758.07361111111, 23758.075, 23758.07638888889, 23758.077777777777, 23758.079166666666, 23758.080555555556, 23758.081944444446, 23758.083333333332, 23758.084722222222, 23758.08611111111, 23758.0875, 23758.088888888888, 23758.090277777777, 23758.091666666667, 23758.093055555557, 23758.094444444443, 23758.095833333333, 23758.097222222223, 23758.098611111112, 23758.1, 23758.10138888889, 23758.102777777778, 23758.104166666668, 23758.105555555554, 23758.106944444444, 23758.108333333334, 23758.109722222223, 23758.11111111111, 23758.1125, 23758.11388888889, 23758.11527777778, 23758.116666666665, 23758.118055555555, 23758.119444444445, 23758.120833333334, 23758.12222222222, 23758.12361111111, 23758.125, 23758.12638888889, 23758.12777777778, 23758.129166666666, 23758.130555555555, 23758.131944444445, 23758.133333333335, 23758.13472222222, 23758.13611111111, 23758.1375, 23758.13888888889, 23758.140277777777, 23758.141666666666, 23758.143055555556, 23758.144444444446, 23758.145833333332, 23758.147222222222, 23758.14861111111, 23758.15, 23758.151388888888, 23758.152777777777, 23758.154166666667, 23758.155555555557, 23758.156944444443, 23758.158333333333, 23758.159722222223, 23758.161111111112, 23758.1625, 23758.16388888889, 23758.165277777778, 23758.166666666668, 23758.168055555554, 23758.169444444444, 23758.170833333334, 23758.172222222223, 23758.17361111111, 23758.175, 23758.17638888889, 23758.17777777778, 23758.179166666665, 23758.180555555555, 23758.181944444445, 23758.183333333334, 23758.18472222222, 23758.18611111111, 23758.1875, 23758.18888888889, 23758.19027777778, 23758.191666666666, 23758.193055555555, 23758.194444444445, 23758.195833333335, 23758.19722222222, 23758.19861111111, 23758.2, 23758.20138888889, 23758.202777777777, 23758.204166666666, 23758.205555555556, 23758.206944444446, 23758.208333333332, 23758.209722222222, 23758.21111111111, 23758.2125, 23758.213888888888, 23758.215277777777, 23758.216666666667, 23758.218055555557, 23758.219444444443, 23758.220833333333, 23758.222222222223, 23758.223611111112, 23758.225, 23758.22638888889, 23758.227777777778, 23758.229166666668, 23758.230555555554, 23758.231944444444, 23758.233333333334, 23758.234722222223, 23758.23611111111, 23758.2375, 23758.23888888889, 23758.24027777778, 23758.241666666665, 23758.243055555555, 23758.244444444445, 23758.245833333334, 23758.24722222222, 23758.24861111111, 23758.25, 23758.25138888889, 23758.25277777778, 23758.254166666666, 23758.255555555555, 23758.256944444445, 23758.258333333335, 23758.25972222222, 23758.26111111111, 23758.2625, 23758.26388888889, 23758.265277777777, 23758.266666666666, 23758.268055555556, 23758.269444444446, 23758.270833333332, 23758.272222222222, 23758.27361111111, 23758.275, 23758.276388888888, 23758.277777777777, 23758.279166666667, 23758.280555555557, 23758.281944444443, 23758.283333333333, 23758.284722222223, 23758.286111111112, 23758.2875, 23758.28888888889, 23758.290277777778, 23758.291666666668, 23758.293055555554, 23758.294444444444, 23758.295833333334, 23758.297222222223, 23758.29861111111, 23758.3, 23758.30138888889, 23758.30277777778, 23758.304166666665, 23758.305555555555, 23758.306944444445, 23758.308333333334, 23758.30972222222, 23758.31111111111, 23758.3125, 23758.31388888889, 23758.31527777778, 23758.316666666666, 23758.318055555555, 23758.319444444445, 23758.320833333335, 23758.32222222222, 23758.32361111111, 23758.325, 23758.32638888889, 23758.327777777777, 23758.329166666666, 23758.330555555556, 23758.331944444446, 23758.333333333332, 23758.334722222222, 23758.33611111111, 23758.3375, 23758.338888888888, 23758.340277777777, 23758.341666666667, 23758.343055555557, 23758.344444444443, 23758.345833333333, 23758.347222222223, 23758.348611111112, 23758.35, 23758.35138888889, 23758.352777777778, 23758.354166666668, 23758.355555555554, 23758.356944444444, 23758.358333333334, 23758.359722222223, 23758.36111111111, 23758.3625, 23758.36388888889, 23758.36527777778, 23758.366666666665, 23758.368055555555, 23758.369444444445, 23758.370833333334, 23758.37222222222, 23758.37361111111, 23758.375, 23758.37638888889, 23758.37777777778, 23758.379166666666, 23758.380555555555, 23758.381944444445, 23758.383333333335, 23758.38472222222, 23758.38611111111, 23758.3875, 23758.38888888889, 23758.390277777777, 23758.391666666666, 23758.393055555556, 23758.394444444446, 23758.395833333332, 23758.397222222222, 23758.39861111111, 23758.4, 23758.401388888888, 23758.402777777777, 23758.404166666667, 23758.405555555557, 23758.406944444443, 23758.408333333333, 23758.409722222223, 23758.411111111112, 23758.4125, 23758.41388888889, 23758.415277777778, 23758.416666666668, 23758.418055555554, 23758.419444444444, 23758.420833333334, 23758.422222222223, 23758.42361111111, 23758.425, 23758.42638888889, 23758.42777777778, 23758.429166666665, 23758.430555555555, 23758.431944444445, 23758.433333333334, 23758.43472222222, 23758.43611111111, 23758.4375, 23758.43888888889, 23758.44027777778, 23758.441666666666, 23758.443055555555, 23758.444444444445, 23758.445833333335, 23758.44722222222, 23758.44861111111, 23758.45, 23758.45138888889, 23758.452777777777, 23758.454166666666, 23758.455555555556, 23758.456944444446, 23758.458333333332, 23758.459722222222, 23758.46111111111, 23758.4625, 23758.463888888888, 23758.465277777777, 23758.466666666667, 23758.468055555557, 23758.469444444443, 23758.470833333333, 23758.472222222223, 23758.473611111112, 23758.475, 23758.47638888889, 23758.477777777778, 23758.479166666668, 23758.480555555554, 23758.481944444444, 23758.483333333334, 23758.484722222223, 23758.48611111111, 23758.4875, 23758.48888888889, 23758.49027777778, 23758.491666666665, 23758.493055555555, 23758.494444444445, 23758.495833333334, 23758.49722222222, 23758.49861111111, 23758.5, 23758.50138888889, 23758.50277777778, 23758.504166666666, 23758.505555555555, 23758.506944444445, 23758.508333333335, 23758.50972222222, 23758.51111111111, 23758.5125, 23758.51388888889, 23758.515277777777, 23758.516666666666, 23758.518055555556, 23758.519444444446, 23758.520833333332, 23758.522222222222, 23758.52361111111, 23758.525, 23758.526388888888, 23758.527777777777, 23758.529166666667, 23758.530555555557, 23758.531944444443, 23758.533333333333, 23758.534722222223, 23758.536111111112, 23758.5375, 23758.53888888889, 23758.540277777778, 23758.541666666668, 23758.543055555554, 23758.544444444444, 23758.545833333334, 23758.547222222223, 23758.54861111111, 23758.55, 23758.55138888889, 23758.55277777778, 23758.554166666665, 23758.555555555555, 23758.556944444445, 23758.558333333334, 23758.55972222222, 23758.56111111111, 23758.5625, 23758.56388888889, 23758.56527777778, 23758.566666666666, 23758.568055555555, 23758.569444444445, 23758.570833333335, 23758.57222222222, 23758.57361111111, 23758.575, 23758.57638888889, 23758.577777777777, 23758.579166666666, 23758.580555555556, 23758.581944444446, 23758.583333333332, 23758.584722222222, 23758.58611111111, 23758.5875, 23758.588888888888, 23758.590277777777, 23758.591666666667, 23758.593055555557, 23758.594444444443, 23758.595833333333, 23758.597222222223, 23758.598611111112, 23758.6, 23758.60138888889, 23758.602777777778, 23758.604166666668, 23758.605555555554, 23758.606944444444, 23758.608333333334, 23758.609722222223, 23758.61111111111, 23758.6125, 23758.61388888889, 23758.61527777778, 23758.616666666665, 23758.618055555555, 23758.619444444445, 23758.620833333334, 23758.62222222222, 23758.62361111111, 23758.625, 23758.62638888889, 23758.62777777778, 23758.629166666666, 23758.630555555555, 23758.631944444445, 23758.633333333335, 23758.63472222222, 23758.63611111111, 23758.6375, 23758.63888888889, 23758.640277777777, 23758.641666666666, 23758.643055555556, 23758.644444444446, 23758.645833333332, 23758.647222222222, 23758.64861111111, 23758.65, 23758.651388888888, 23758.652777777777, 23758.654166666667, 23758.655555555557, 23758.656944444443, 23758.658333333333, 23758.659722222223, 23758.661111111112, 23758.6625, 23758.66388888889, 23758.665277777778, 23758.666666666668, 23758.668055555554, 23758.669444444444, 23758.670833333334, 23758.672222222223, 23758.67361111111, 23758.675, 23758.67638888889, 23758.67777777778, 23758.679166666665, 23758.680555555555, 23758.681944444445, 23758.683333333334, 23758.68472222222, 23758.68611111111, 23758.6875, 23758.68888888889, 23758.69027777778, 23758.691666666666, 23758.693055555555, 23758.694444444445, 23758.695833333335, 23758.69722222222, 23758.69861111111, 23758.7, 23758.70138888889, 23758.702777777777, 23758.704166666666, 23758.705555555556, 23758.706944444446, 23758.708333333332, 23758.709722222222, 23758.71111111111, 23758.7125, 23758.713888888888, 23758.715277777777, 23758.716666666667, 23758.718055555557, 23758.719444444443, 23758.720833333333, 23758.722222222223, 23758.723611111112, 23758.725, 23758.72638888889, 23758.727777777778, 23758.729166666668, 23758.730555555554, 23758.731944444444, 23758.733333333334, 23758.734722222223, 23758.73611111111, 23758.7375, 23758.73888888889, 23758.74027777778, 23758.741666666665, 23758.743055555555, 23758.744444444445, 23758.745833333334, 23758.74722222222, 23758.74861111111, 23758.75, 23758.75138888889, 23758.75277777778, 23758.754166666666, 23758.755555555555, 23758.756944444445, 23758.758333333335, 23758.75972222222, 23758.76111111111, 23758.7625, 23758.76388888889, 23758.765277777777, 23758.766666666666, 23758.768055555556, 23758.769444444446, 23758.770833333332, 23758.772222222222, 23758.77361111111, 23758.775, 23758.776388888888, 23758.777777777777, 23758.779166666667, 23758.780555555557, 23758.781944444443, 23758.783333333333, 23758.784722222223, 23758.786111111112, 23758.7875, 23758.78888888889, 23758.790277777778, 23758.791666666668, 23758.793055555554, 23758.794444444444, 23758.795833333334, 23758.797222222223, 23758.79861111111, 23758.8, 23758.80138888889, 23758.80277777778, 23758.804166666665, 23758.805555555555, 23758.806944444445, 23758.808333333334, 23758.80972222222, 23758.81111111111, 23758.8125, 23758.81388888889, 23758.81527777778, 23758.816666666666, 23758.818055555555, 23758.819444444445, 23758.820833333335, 23758.82222222222, 23758.82361111111, 23758.825, 23758.82638888889, 23758.827777777777, 23758.829166666666, 23758.830555555556, 23758.831944444446, 23758.833333333332, 23758.834722222222, 23758.83611111111, 23758.8375, 23758.838888888888, 23758.840277777777, 23758.841666666667, 23758.843055555557, 23758.844444444443, 23758.845833333333, 23758.847222222223, 23758.848611111112, 23758.85, 23758.85138888889, 23758.852777777778, 23758.854166666668, 23758.855555555554, 23758.856944444444, 23758.858333333334, 23758.859722222223, 23758.86111111111, 23758.8625, 23758.86388888889, 23758.86527777778, 23758.866666666665, 23758.868055555555, 23758.869444444445, 23758.870833333334, 23758.87222222222, 23758.87361111111, 23758.875, 23758.87638888889, 23758.87777777778, 23758.879166666666, 23758.880555555555, 23758.881944444445, 23758.883333333335, 23758.88472222222, 23758.88611111111, 23758.8875, 23758.88888888889, 23758.890277777777, 23758.891666666666, 23758.893055555556, 23758.894444444446, 23758.895833333332, 23758.897222222222, 23758.89861111111, 23758.9, 23758.901388888888, 23758.902777777777, 23758.904166666667, 23758.905555555557, 23758.906944444443, 23758.908333333333, 23758.909722222223, 23758.911111111112, 23758.9125, 23758.91388888889, 23758.915277777778, 23758.916666666668, 23758.918055555554, 23758.919444444444, 23758.920833333334, 23758.922222222223, 23758.92361111111, 23758.925, 23758.92638888889, 23758.92777777778, 23758.929166666665, 23758.930555555555, 23758.931944444445, 23758.933333333334, 23758.93472222222, 23758.93611111111, 23758.9375, 23758.93888888889, 23758.94027777778, 23758.941666666666, 23758.943055555555, 23758.944444444445, 23758.945833333335, 23758.94722222222, 23758.94861111111, 23758.95, 23758.95138888889, 23758.952777777777, 23758.954166666666, 23758.955555555556, 23758.956944444446, 23758.958333333332, 23758.959722222222, 23758.96111111111, 23758.9625, 23758.963888888888, 23758.965277777777, 23758.966666666667, 23758.968055555557, 23758.969444444443, 23758.970833333333, 23758.972222222223, 23758.973611111112, 23758.975, 23758.97638888889, 23758.977777777778, 23758.979166666668, 23758.980555555554, 23758.981944444444, 23758.983333333334, 23758.984722222223, 23758.98611111111, 23758.9875, 23758.98888888889, 23758.99027777778, 23758.991666666665, 23758.993055555555, 23758.994444444445, 23758.995833333334, 23758.99722222222, 23758.99861111111, 23759.0, 23759.00138888889, 23759.00277777778, 23759.004166666666, 23759.005555555555, 23759.006944444445, 23759.008333333335, 23759.00972222222, 23759.01111111111, 23759.0125, 23759.01388888889, 23759.015277777777, 23759.016666666666, 23759.018055555556, 23759.019444444446, 23759.020833333332, 23759.022222222222, 23759.02361111111, 23759.025, 23759.026388888888, 23759.027777777777, 23759.029166666667, 23759.030555555557, 23759.031944444443, 23759.033333333333, 23759.034722222223, 23759.036111111112, 23759.0375, 23759.03888888889, 23759.040277777778, 23759.041666666668, 23759.043055555554, 23759.044444444444, 23759.045833333334, 23759.047222222223, 23759.04861111111, 23759.05, 23759.05138888889, 23759.05277777778, 23759.054166666665, 23759.055555555555, 23759.056944444445, 23759.058333333334, 23759.05972222222, 23759.06111111111, 23759.0625, 23759.06388888889, 23759.06527777778, 23759.066666666666, 23759.068055555555, 23759.069444444445, 23759.070833333335, 23759.07222222222, 23759.07361111111, 23759.075, 23759.07638888889, 23759.077777777777, 23759.079166666666, 23759.080555555556, 23759.081944444446, 23759.083333333332, 23759.084722222222, 23759.08611111111, 23759.0875, 23759.088888888888, 23759.090277777777, 23759.091666666667, 23759.093055555557, 23759.094444444443, 23759.095833333333, 23759.097222222223, 23759.098611111112, 23759.1, 23759.10138888889, 23759.102777777778, 23759.104166666668, 23759.105555555554, 23759.106944444444, 23759.108333333334, 23759.109722222223, 23759.11111111111, 23759.1125, 23759.11388888889, 23759.11527777778, 23759.116666666665, 23759.118055555555, 23759.119444444445, 23759.120833333334, 23759.12222222222, 23759.12361111111, 23759.125, 23759.12638888889, 23759.12777777778, 23759.129166666666, 23759.130555555555, 23759.131944444445, 23759.133333333335, 23759.13472222222, 23759.13611111111, 23759.1375, 23759.13888888889, 23759.140277777777, 23759.141666666666, 23759.143055555556, 23759.144444444446, 23759.145833333332, 23759.147222222222, 23759.14861111111, 23759.15, 23759.151388888888, 23759.152777777777, 23759.154166666667, 23759.155555555557, 23759.156944444443, 23759.158333333333, 23759.159722222223, 23759.161111111112, 23759.1625, 23759.16388888889, 23759.165277777778, 23759.166666666668, 23759.168055555554, 23759.169444444444, 23759.170833333334, 23759.172222222223, 23759.17361111111, 23759.175, 23759.17638888889, 23759.17777777778, 23759.179166666665, 23759.180555555555, 23759.181944444445, 23759.183333333334, 23759.18472222222, 23759.18611111111, 23759.1875, 23759.18888888889, 23759.19027777778, 23759.191666666666, 23759.193055555555, 23759.194444444445, 23759.195833333335, 23759.19722222222, 23759.19861111111, 23759.2, 23759.20138888889, 23759.202777777777, 23759.204166666666, 23759.205555555556, 23759.206944444446, 23759.208333333332, 23759.209722222222, 23759.21111111111, 23759.2125, 23759.213888888888, 23759.215277777777, 23759.216666666667, 23759.218055555557, 23759.219444444443, 23759.220833333333, 23759.222222222223, 23759.223611111112, 23759.225, 23759.22638888889, 23759.227777777778, 23759.229166666668, 23759.230555555554, 23759.231944444444, 23759.233333333334, 23759.234722222223, 23759.23611111111, 23759.2375, 23759.23888888889, 23759.24027777778, 23759.241666666665, 23759.243055555555, 23759.244444444445, 23759.245833333334, 23759.24722222222, 23759.24861111111, 23759.25, 23759.25138888889, 23759.25277777778, 23759.254166666666, 23759.255555555555, 23759.256944444445, 23759.258333333335, 23759.25972222222, 23759.26111111111, 23759.2625, 23759.26388888889, 23759.265277777777, 23759.266666666666, 23759.268055555556, 23759.269444444446, 23759.270833333332, 23759.272222222222, 23759.27361111111, 23759.275, 23759.276388888888, 23759.277777777777, 23759.279166666667, 23759.280555555557, 23759.281944444443, 23759.283333333333, 23759.284722222223, 23759.286111111112, 23759.2875, 23759.28888888889, 23759.290277777778, 23759.291666666668, 23759.293055555554, 23759.294444444444, 23759.295833333334, 23759.297222222223, 23759.29861111111, 23759.3, 23759.30138888889, 23759.30277777778, 23759.304166666665, 23759.305555555555, 23759.306944444445, 23759.308333333334, 23759.30972222222, 23759.31111111111, 23759.3125, 23759.31388888889, 23759.31527777778, 23759.316666666666, 23759.318055555555, 23759.319444444445, 23759.320833333335, 23759.32222222222, 23759.32361111111, 23759.325, 23759.32638888889, 23759.327777777777, 23759.329166666666, 23759.330555555556, 23759.331944444446, 23759.333333333332, 23759.334722222222, 23759.33611111111, 23759.3375, 23759.338888888888, 23759.340277777777, 23759.341666666667, 23759.343055555557, 23759.344444444443, 23759.345833333333, 23759.347222222223, 23759.348611111112, 23759.35, 23759.35138888889, 23759.352777777778, 23759.354166666668, 23759.355555555554, 23759.356944444444, 23759.358333333334, 23759.359722222223, 23759.36111111111, 23759.3625, 23759.36388888889, 23759.36527777778, 23759.366666666665, 23759.368055555555, 23759.369444444445, 23759.370833333334, 23759.37222222222, 23759.37361111111, 23759.375, 23759.37638888889, 23759.37777777778, 23759.379166666666, 23759.380555555555, 23759.381944444445, 23759.383333333335, 23759.38472222222, 23759.38611111111, 23759.3875, 23759.38888888889, 23759.390277777777, 23759.391666666666, 23759.393055555556, 23759.394444444446, 23759.395833333332, 23759.397222222222, 23759.39861111111, 23759.4, 23759.401388888888, 23759.402777777777, 23759.404166666667, 23759.405555555557, 23759.406944444443, 23759.408333333333, 23759.409722222223, 23759.411111111112, 23759.4125, 23759.41388888889, 23759.415277777778, 23759.416666666668, 23759.418055555554, 23759.419444444444, 23759.420833333334, 23759.422222222223, 23759.42361111111, 23759.425, 23759.42638888889, 23759.42777777778, 23759.429166666665, 23759.430555555555, 23759.431944444445, 23759.433333333334, 23759.43472222222, 23759.43611111111, 23759.4375, 23759.43888888889, 23759.44027777778, 23759.441666666666, 23759.443055555555, 23759.444444444445, 23759.445833333335, 23759.44722222222, 23759.44861111111, 23759.45, 23759.45138888889, 23759.452777777777, 23759.454166666666, 23759.455555555556, 23759.456944444446, 23759.458333333332, 23759.459722222222, 23759.46111111111, 23759.4625, 23759.463888888888, 23759.465277777777, 23759.466666666667, 23759.468055555557, 23759.469444444443, 23759.470833333333, 23759.472222222223, 23759.473611111112, 23759.475, 23759.47638888889, 23759.477777777778, 23759.479166666668, 23759.480555555554, 23759.481944444444, 23759.483333333334, 23759.484722222223, 23759.48611111111, 23759.4875, 23759.48888888889, 23759.49027777778, 23759.491666666665, 23759.493055555555, 23759.494444444445, 23759.495833333334, 23759.49722222222, 23759.49861111111, 23759.5, 23759.50138888889, 23759.50277777778, 23759.504166666666, 23759.505555555555, 23759.506944444445, 23759.508333333335, 23759.50972222222, 23759.51111111111, 23759.5125, 23759.51388888889, 23759.515277777777, 23759.516666666666, 23759.518055555556, 23759.519444444446, 23759.520833333332, 23759.522222222222, 23759.52361111111, 23759.525, 23759.526388888888, 23759.527777777777, 23759.529166666667, 23759.530555555557, 23759.531944444443, 23759.533333333333, 23759.534722222223, 23759.536111111112, 23759.5375, 23759.53888888889, 23759.540277777778, 23759.541666666668, 23759.543055555554, 23759.544444444444, 23759.545833333334, 23759.547222222223, 23759.54861111111, 23759.55, 23759.55138888889, 23759.55277777778, 23759.554166666665, 23759.555555555555, 23759.556944444445, 23759.558333333334, 23759.55972222222, 23759.56111111111, 23759.5625, 23759.56388888889, 23759.56527777778, 23759.566666666666, 23759.568055555555, 23759.569444444445, 23759.570833333335, 23759.57222222222, 23759.57361111111, 23759.575, 23759.57638888889, 23759.577777777777, 23759.579166666666, 23759.580555555556, 23759.581944444446, 23759.583333333332, 23759.584722222222, 23759.58611111111, 23759.5875, 23759.588888888888, 23759.590277777777, 23759.591666666667, 23759.593055555557, 23759.594444444443, 23759.595833333333, 23759.597222222223, 23759.598611111112, 23759.6, 23759.60138888889, 23759.602777777778, 23759.604166666668, 23759.605555555554, 23759.606944444444, 23759.608333333334, 23759.609722222223, 23759.61111111111, 23759.6125, 23759.61388888889, 23759.61527777778, 23759.616666666665, 23759.618055555555, 23759.619444444445, 23759.620833333334, 23759.62222222222, 23759.62361111111, 23759.625, 23759.62638888889, 23759.62777777778, 23759.629166666666, 23759.630555555555, 23759.631944444445, 23759.633333333335, 23759.63472222222, 23759.63611111111, 23759.6375, 23759.63888888889, 23759.640277777777, 23759.641666666666, 23759.643055555556, 23759.644444444446, 23759.645833333332, 23759.647222222222, 23759.64861111111, 23759.65, 23759.651388888888, 23759.652777777777, 23759.654166666667, 23759.655555555557, 23759.656944444443, 23759.658333333333, 23759.659722222223, 23759.661111111112, 23759.6625, 23759.66388888889, 23759.665277777778, 23759.666666666668, 23759.668055555554, 23759.669444444444, 23759.670833333334, 23759.672222222223, 23759.67361111111, 23759.675, 23759.67638888889, 23759.67777777778, 23759.679166666665, 23759.680555555555, 23759.681944444445, 23759.683333333334, 23759.68472222222, 23759.68611111111, 23759.6875, 23759.68888888889, 23759.69027777778, 23759.691666666666, 23759.693055555555, 23759.694444444445, 23759.695833333335, 23759.69722222222, 23759.69861111111, 23759.7, 23759.70138888889, 23759.702777777777, 23759.704166666666, 23759.705555555556, 23759.706944444446, 23759.708333333332, 23759.709722222222, 23759.71111111111, 23759.7125, 23759.713888888888, 23759.715277777777, 23759.716666666667, 23759.718055555557, 23759.719444444443, 23759.720833333333, 23759.722222222223, 23759.723611111112, 23759.725, 23759.72638888889, 23759.727777777778, 23759.729166666668, 23759.730555555554, 23759.731944444444, 23759.733333333334, 23759.734722222223, 23759.73611111111, 23759.7375, 23759.73888888889, 23759.74027777778, 23759.741666666665, 23759.743055555555, 23759.744444444445, 23759.745833333334, 23759.74722222222, 23759.74861111111, 23759.75, 23759.75138888889, 23759.75277777778, 23759.754166666666, 23759.755555555555, 23759.756944444445, 23759.758333333335, 23759.75972222222, 23759.76111111111, 23759.7625, 23759.76388888889, 23759.765277777777, 23759.766666666666, 23759.768055555556, 23759.769444444446, 23759.770833333332, 23759.772222222222, 23759.77361111111, 23759.775, 23759.776388888888, 23759.777777777777, 23759.779166666667, 23759.780555555557, 23759.781944444443, 23759.783333333333, 23759.784722222223, 23759.786111111112, 23759.7875, 23759.78888888889, 23759.790277777778, 23759.791666666668, 23759.793055555554, 23759.794444444444, 23759.795833333334, 23759.797222222223, 23759.79861111111, 23759.8, 23759.80138888889, 23759.80277777778, 23759.804166666665, 23759.805555555555, 23759.806944444445, 23759.808333333334, 23759.80972222222, 23759.81111111111, 23759.8125, 23759.81388888889, 23759.81527777778, 23759.816666666666, 23759.818055555555, 23759.819444444445, 23759.820833333335, 23759.82222222222, 23759.82361111111, 23759.825, 23759.82638888889, 23759.827777777777, 23759.829166666666, 23759.830555555556, 23759.831944444446, 23759.833333333332, 23759.834722222222, 23759.83611111111, 23759.8375, 23759.838888888888, 23759.840277777777, 23759.841666666667, 23759.843055555557, 23759.844444444443, 23759.845833333333, 23759.847222222223, 23759.848611111112, 23759.85, 23759.85138888889, 23759.852777777778, 23759.854166666668, 23759.855555555554, 23759.856944444444, 23759.858333333334, 23759.859722222223, 23759.86111111111, 23759.8625, 23759.86388888889, 23759.86527777778, 23759.866666666665, 23759.868055555555, 23759.869444444445, 23759.870833333334, 23759.87222222222, 23759.87361111111, 23759.875, 23759.87638888889, 23759.87777777778, 23759.879166666666, 23759.880555555555, 23759.881944444445, 23759.883333333335, 23759.88472222222, 23759.88611111111, 23759.8875, 23759.88888888889, 23759.890277777777, 23759.891666666666, 23759.893055555556, 23759.894444444446, 23759.895833333332, 23759.897222222222, 23759.89861111111, 23759.9, 23759.901388888888, 23759.902777777777, 23759.904166666667, 23759.905555555557, 23759.906944444443, 23759.908333333333, 23759.909722222223, 23759.911111111112, 23759.9125, 23759.91388888889, 23759.915277777778, 23759.916666666668, 23759.918055555554, 23759.919444444444, 23759.920833333334, 23759.922222222223, 23759.92361111111, 23759.925, 23759.92638888889, 23759.92777777778, 23759.929166666665, 23759.930555555555, 23759.931944444445, 23759.933333333334, 23759.93472222222, 23759.93611111111, 23759.9375, 23759.93888888889, 23759.94027777778, 23759.941666666666, 23759.943055555555, 23759.944444444445, 23759.945833333335, 23759.94722222222, 23759.94861111111, 23759.95, 23759.95138888889, 23759.952777777777, 23759.954166666666, 23759.955555555556, 23759.956944444446, 23759.958333333332, 23759.959722222222, 23759.96111111111, 23759.9625, 23759.963888888888, 23759.965277777777, 23759.966666666667, 23759.968055555557, 23759.969444444443, 23759.970833333333, 23759.972222222223, 23759.973611111112, 23759.975, 23759.97638888889, 23759.977777777778, 23759.979166666668, 23759.980555555554, 23759.981944444444, 23759.983333333334, 23759.984722222223, 23759.98611111111, 23759.9875, 23759.98888888889, 23759.99027777778, 23759.991666666665, 23759.993055555555, 23759.994444444445, 23759.995833333334, 23759.99722222222, 23759.99861111111, 23760.0, 23760.00138888889, 23760.00277777778, 23760.004166666666, 23760.005555555555, 23760.006944444445, 23760.008333333335, 23760.00972222222, 23760.01111111111, 23760.0125, 23760.01388888889, 23760.015277777777, 23760.016666666666, 23760.018055555556, 23760.019444444446, 23760.020833333332, 23760.022222222222, 23760.02361111111, 23760.025, 23760.026388888888, 23760.027777777777, 23760.029166666667, 23760.030555555557, 23760.031944444443, 23760.033333333333, 23760.034722222223, 23760.036111111112, 23760.0375, 23760.03888888889, 23760.040277777778, 23760.041666666668, 23760.043055555554, 23760.044444444444, 23760.045833333334, 23760.047222222223, 23760.04861111111, 23760.05, 23760.05138888889, 23760.05277777778, 23760.054166666665, 23760.055555555555, 23760.056944444445, 23760.058333333334, 23760.05972222222, 23760.06111111111, 23760.0625, 23760.06388888889, 23760.06527777778, 23760.066666666666, 23760.068055555555, 23760.069444444445, 23760.070833333335, 23760.07222222222, 23760.07361111111, 23760.075, 23760.07638888889, 23760.077777777777, 23760.079166666666, 23760.080555555556, 23760.081944444446, 23760.083333333332, 23760.084722222222, 23760.08611111111, 23760.0875, 23760.088888888888, 23760.090277777777, 23760.091666666667, 23760.093055555557, 23760.094444444443, 23760.095833333333, 23760.097222222223, 23760.098611111112, 23760.1, 23760.10138888889, 23760.102777777778, 23760.104166666668, 23760.105555555554, 23760.106944444444, 23760.108333333334, 23760.109722222223, 23760.11111111111, 23760.1125, 23760.11388888889, 23760.11527777778, 23760.116666666665, 23760.118055555555, 23760.119444444445, 23760.120833333334, 23760.12222222222, 23760.12361111111, 23760.125, 23760.12638888889, 23760.12777777778, 23760.129166666666, 23760.130555555555, 23760.131944444445, 23760.133333333335, 23760.13472222222, 23760.13611111111, 23760.1375, 23760.13888888889, 23760.140277777777, 23760.141666666666, 23760.143055555556, 23760.144444444446, 23760.145833333332, 23760.147222222222, 23760.14861111111, 23760.15, 23760.151388888888, 23760.152777777777, 23760.154166666667, 23760.155555555557, 23760.156944444443, 23760.158333333333, 23760.159722222223, 23760.161111111112, 23760.1625, 23760.16388888889, 23760.165277777778, 23760.166666666668, 23760.168055555554, 23760.169444444444, 23760.170833333334, 23760.172222222223, 23760.17361111111, 23760.175, 23760.17638888889, 23760.17777777778, 23760.179166666665, 23760.180555555555, 23760.181944444445, 23760.183333333334, 23760.18472222222, 23760.18611111111, 23760.1875, 23760.18888888889, 23760.19027777778, 23760.191666666666, 23760.193055555555, 23760.194444444445, 23760.195833333335, 23760.19722222222, 23760.19861111111, 23760.2, 23760.20138888889, 23760.202777777777, 23760.204166666666, 23760.205555555556, 23760.206944444446, 23760.208333333332, 23760.209722222222, 23760.21111111111, 23760.2125, 23760.213888888888, 23760.215277777777, 23760.216666666667, 23760.218055555557, 23760.219444444443, 23760.220833333333, 23760.222222222223, 23760.223611111112, 23760.225, 23760.22638888889, 23760.227777777778, 23760.229166666668, 23760.230555555554, 23760.231944444444, 23760.233333333334, 23760.234722222223, 23760.23611111111, 23760.2375, 23760.23888888889, 23760.24027777778, 23760.241666666665, 23760.243055555555, 23760.244444444445, 23760.245833333334, 23760.24722222222, 23760.24861111111, 23760.25, 23760.25138888889, 23760.25277777778, 23760.254166666666, 23760.255555555555, 23760.256944444445, 23760.258333333335, 23760.25972222222, 23760.26111111111, 23760.2625, 23760.26388888889, 23760.265277777777, 23760.266666666666, 23760.268055555556, 23760.269444444446, 23760.270833333332, 23760.272222222222, 23760.27361111111, 23760.275, 23760.276388888888, 23760.277777777777, 23760.279166666667, 23760.280555555557, 23760.281944444443, 23760.283333333333, 23760.284722222223, 23760.286111111112, 23760.2875, 23760.28888888889, 23760.290277777778, 23760.291666666668, 23760.293055555554, 23760.294444444444, 23760.295833333334, 23760.297222222223, 23760.29861111111, 23760.3, 23760.30138888889, 23760.30277777778}
LATITUDE =-31.7285666667
LONGITUDE =115.0371
NOMINAL_DEPTH =196.0
TEMP =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
TEMP_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
CNDC =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
CNDC_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PSAL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PSAL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
PRES =
  {218.4761, 218.4889, 218.4929, 218.4937, 218.494, 218.4986, 218.4982, 218.5084, 218.5045, 218.5, 218.4894, 218.5053, 218.4765, 218.4832, 218.4905, 218.4991, 218.4958, 218.4993, 218.4989, 218.5014, 218.4905, 218.4987, 218.4944, 218.4904, 218.4943, 218.4847, 218.4894, 218.4836, 218.4851, 218.4901, 218.5081, 218.5071, 218.5058, 218.503, 218.5173, 218.5014, 218.5097, 218.5125, 218.5156, 218.5112, 218.4996, 218.512, 218.5118, 218.5133, 218.5152, 218.5132, 218.5268, 218.5234, 218.5206, 218.5245, 218.538, 218.556, 218.5223, 218.5389, 218.5354, 218.542, 218.5284, 218.539, 218.5501, 218.54, 218.5503, 218.5397, 218.5637, 218.558, 218.5394, 218.5587, 218.549, 218.566, 218.5664, 218.5585, 218.5684, 218.5794, 218.5755, 218.5755, 218.5629, 218.5795, 218.5636, 218.5981, 218.5778, 218.5762, 218.5904, 218.5737, 218.577, 218.5914, 218.5802, 218.5872, 218.5831, 218.5831, 218.5741, 218.5744, 218.5966, 218.5836, 218.5932, 218.5951, 218.5884, 218.6028, 218.6119, 218.6045, 218.6183, 218.592, 218.6128, 218.6133, 218.6036, 218.6114, 218.6061, 218.6031, 218.6233, 218.6033, 218.6051, 218.6183, 218.5929, 218.6106, 218.6149, 218.6215, 218.6165, 218.6053, 218.6165, 218.6141, 218.624, 218.6144, 218.6262, 218.6292, 218.6499, 218.6287, 218.6306, 218.6296, 218.6317, 218.6272, 218.6218, 218.639, 218.6346, 218.6359, 218.6454, 218.64, 218.6375, 218.644, 218.6464, 218.6353, 218.6425, 218.6362, 218.6353, 218.6546, 218.6542, 218.6635, 218.6386, 218.6457, 218.6572, 218.6413, 218.6431, 218.6403, 218.6586, 218.6713, 218.6504, 218.6444, 218.6516, 218.6718, 218.6737, 218.6697, 218.6802, 218.6721, 218.6646, 218.6707, 218.6709, 218.6628, 218.672, 218.6764, 218.6868, 218.6749, 218.6734, 218.6738, 218.7044, 218.6765, 218.6711, 218.6788, 218.6776, 218.6847, 218.6871, 218.6835, 218.7007, 218.6954, 218.6778, 218.6834, 218.6787, 218.6859, 218.686, 218.6726, 218.6929, 218.6928, 218.6938, 218.6928, 218.7009, 218.6801, 218.6819, 218.6845, 218.7104, 218.6886, 218.7047, 218.702, 218.7089, 218.7091, 218.6997, 218.7037, 218.712, 218.7092, 218.721, 218.7201, 218.7105, 218.6978, 218.7306, 218.6976, 218.7006, 218.7069, 218.7139, 218.7154, 218.7179, 218.7277, 218.7101, 218.7067, 218.7184, 218.7083, 218.7255, 218.7297, 218.7201, 218.7182, 218.7232, 218.716, 218.719, 218.71, 218.7326, 218.7242, 218.7303, 218.7204, 218.7298, 218.7331, 218.7265, 218.7234, 218.7389, 218.7534, 218.7216, 218.7333, 218.7234, 218.7441, 218.7377, 218.7573, 218.7309, 218.7397, 218.7446, 218.7433, 218.7349, 218.748, 218.7578, 218.7595, 218.7289, 218.7537, 218.757, 218.7595, 218.7709, 218.7528, 218.7706, 218.7604, 218.772, 218.7542, 218.7567, 218.7615, 218.7642, 218.7544, 218.7677, 218.7763, 218.7667, 218.7766, 218.7864, 218.7731, 218.7723, 218.7713, 218.7859, 218.7782, 218.7807, 218.7501, 218.7746, 218.776, 218.7804, 218.7681, 218.7749, 218.7808, 218.7708, 218.7851, 218.7867, 218.7808, 218.7802, 218.7813, 218.7721, 218.7942, 218.8008, 218.7988, 218.7934, 218.7929, 218.783, 218.7791, 218.7928, 218.7783, 218.7895, 218.7977, 218.7656, 218.7858, 218.7904, 218.7729, 218.7975, 218.7772, 218.8024, 218.7925, 218.7909, 218.7914, 218.7812, 218.7796, 218.7864, 218.7855, 218.7935, 218.7896, 218.7695, 218.7985, 218.7791, 218.794, 218.7919, 218.7866, 218.7949, 218.8055, 218.7904, 218.7813, 218.7902, 218.7912, 218.7931, 218.7829, 218.7743, 218.7869, 218.7856, 218.7906, 218.7876, 218.788, 218.7789, 218.7849, 218.7803, 218.7708, 218.7801, 218.7959, 218.7645, 218.7911, 218.7864, 218.7966, 218.7689, 218.7918, 218.7899, 218.7895, 218.7795, 218.7862, 218.8005, 218.7731, 218.7863, 218.7754, 218.7873, 218.7999, 218.7816, 218.7858, 218.7938, 218.7811, 218.7887, 218.7814, 218.7915, 218.7905, 218.7773, 218.782, 218.7839, 218.774, 218.7798, 218.7786, 218.776, 218.7647, 218.7692, 218.7675, 218.7591, 218.766, 218.7607, 218.7733, 218.7707, 218.7704, 218.7579, 218.7529, 218.7691, 218.7496, 218.7553, 218.7622, 218.7564, 218.753, 218.7656, 218.7442, 218.7617, 218.7668, 218.7434, 218.745, 218.7525, 218.7443, 218.7289, 218.7362, 218.7375, 218.7509, 218.7348, 218.7355, 218.7457, 218.7256, 218.7319, 218.7405, 218.7328, 218.7223, 218.7357, 218.7298, 218.7305, 218.7135, 218.7311, 218.7192, 218.7171, 218.7206, 218.7179, 218.7116, 218.7025, 218.7251, 218.7145, 218.7154, 218.7042, 218.6914, 218.7082, 218.6972, 218.6988, 218.6955, 218.7014, 218.6954, 218.6928, 218.6844, 218.6888, 218.6856, 218.7004, 218.6886, 218.6753, 218.6899, 218.6843, 218.6866, 218.6812, 218.6809, 218.6739, 218.6623, 218.6813, 218.6723, 218.6729, 218.6679, 218.6515, 218.6539, 218.6635, 218.6736, 218.6447, 218.6488, 218.6588, 218.6466, 218.6467, 218.6517, 218.6572, 218.6498, 218.6428, 218.6387, 218.6436, 218.639, 218.6455, 218.6219, 218.6303, 218.6376, 218.6301, 218.6164, 218.6302, 218.6177, 218.6271, 218.6225, 218.6127, 218.6284, 218.6145, 218.6337, 218.6027, 218.617, 218.6156, 218.6179, 218.6056, 218.5989, 218.607, 218.5947, 218.5914, 218.6062, 218.588, 218.5942, 218.58, 218.5806, 218.5988, 218.5844, 218.5864, 218.59, 218.5595, 218.5994, 218.5844, 218.5871, 218.5729, 218.5843, 218.5807, 218.568, 218.5798, 218.5793, 218.5806, 218.5585, 218.5791, 218.5633, 218.574, 218.5785, 218.559, 218.5401, 218.5629, 218.5573, 218.5519, 218.5457, 218.5761, 218.5578, 218.5507, 218.5489, 218.5523, 218.5497, 218.5504, 218.544, 218.5447, 218.5326, 218.5428, 218.5308, 218.5485, 218.526, 218.5455, 218.5427, 218.5351, 218.5385, 218.5444, 218.5435, 218.5406, 218.5222, 218.5166, 218.5322, 218.5271, 218.5259, 218.5279, 218.5131, 218.5255, 218.5219, 218.5199, 218.5149, 218.5314, 218.5212, 218.515, 218.5134, 218.5092, 218.5168, 218.4986, 218.5165, 218.4978, 218.503, 218.515, 218.4892, 218.5001, 218.5084, 218.5053, 218.4908, 218.5099, 218.4809, 218.4959, 218.4948, 218.499, 218.476, 218.4747, 218.4828, 218.4827, 218.4876, 218.4677, 218.4819, 218.4902, 218.4634, 218.4782, 218.4691, 218.503, 218.4515, 218.4621, 218.478, 218.4737, 218.4594, 218.479, 218.4513, 218.4668, 218.4798, 218.4628, 218.4732, 218.4715, 218.4685, 218.4705, 218.4581, 218.4637, 218.4573, 218.4576, 218.4635, 218.4599, 218.4474, 218.4386, 218.4474, 218.447, 218.4536, 218.4304, 218.4371, 218.4315, 218.4374, 218.4496, 218.4425, 218.4443, 218.4438, 218.4311, 218.4286, 218.437, 218.4413, 218.4404, 218.4297, 218.435, 218.4277, 218.4224, 218.4368, 218.4275, 218.4452, 218.4398, 218.4421, 218.4342, 218.4179, 218.4209, 218.4194, 218.4407, 218.4291, 218.4278, 218.4207, 218.4216, 218.4337, 218.4361, 218.4326, 218.4264, 218.4336, 218.4277, 218.4209, 218.424, 218.4311, 218.4314, 218.4177, 218.4292, 218.4292, 218.4195, 218.4148, 218.4348, 218.4362, 218.4351, 218.4317, 218.4269, 218.4204, 218.4324, 218.4248, 218.4263, 218.4143, 218.4146, 218.419, 218.4444, 218.4241, 218.4458, 218.4266, 218.4436, 218.433, 218.4218, 218.4345, 218.4435, 218.436, 218.4456, 218.4526, 218.4533, 218.4374, 218.4512, 218.4427, 218.4508, 218.4503, 218.4566, 218.4508, 218.4519, 218.4539, 218.4443, 218.4428, 218.458, 218.4463, 218.4584, 218.4435, 218.4604, 218.476, 218.4595, 218.4652, 218.4483, 218.4433, 218.4537, 218.4426, 218.4513, 218.4544, 218.4448, 218.454, 218.4465, 218.4452, 218.4523, 218.4489, 218.4616, 218.4509, 218.4508, 218.4581, 218.4499, 218.4563, 218.4626, 218.4699, 218.4442, 218.4548, 218.4688, 218.4753, 218.4675, 218.4506, 218.4713, 218.4641, 218.477, 218.4662, 218.4624, 218.4782, 218.4788, 218.4797, 218.4842, 218.4706, 218.4612, 218.4772, 218.4858, 218.495, 218.4854, 218.4776, 218.4875, 218.4725, 218.4836, 218.4813, 218.486, 218.4966, 218.4887, 218.4957, 218.4858, 218.487, 218.5018, 218.5204, 218.4923, 218.5004, 218.5046, 218.4901, 218.4963, 218.4929, 218.5075, 218.4924, 218.5073, 218.4944, 218.5018, 218.5023, 218.5051, 218.4981, 218.4908, 218.4928, 218.5169, 218.5046, 218.5049, 218.5116, 218.5137, 218.5048, 218.5061, 218.5175, 218.5322, 218.5331, 218.5286, 218.5134, 218.5093, 218.5275, 218.5187, 218.5205, 218.5235, 218.5435, 218.5256, 218.5131, 218.5238, 218.5199, 218.5345, 218.5239, 218.5159, 218.5359, 218.5225, 218.525, 218.5468, 218.5336, 218.531, 218.5304, 218.541, 218.551, 218.5474, 218.5434, 218.5542, 218.5494, 218.5561, 218.5634, 218.5505, 218.5506, 218.5614, 218.5617, 218.5678, 218.5688, 218.5625, 218.5519, 218.5598, 218.5701, 218.5719, 218.5501, 218.5686, 218.5843, 218.5675, 218.5646, 218.5768, 218.5882, 218.5664, 218.5815, 218.5745, 218.5804, 218.591, 218.5684, 218.5683, 218.5895, 218.5908, 218.5886, 218.5851, 218.5872, 218.5932, 218.5851, 218.5771, 218.5991, 218.5834, 218.6015, 218.5896, 218.5882, 218.596, 218.5806, 218.5968, 218.6106, 218.6143, 218.6011, 218.5981, 218.6125, 218.6263, 218.6169, 218.6325, 218.6103, 218.6183, 218.6123, 218.6107, 218.6191, 218.6317, 218.6308, 218.6178, 218.6369, 218.6073, 218.6227, 218.627, 218.6366, 218.6425, 218.6304, 218.6212, 218.6346, 218.6435, 218.6241, 218.6219, 218.6318, 218.6196, 218.6526, 218.6391, 218.6428, 218.6488, 218.648, 218.6483, 218.6487, 218.6473, 218.6644, 218.6414, 218.6511, 218.6615, 218.6461, 218.6677, 218.6629, 218.677, 218.6777, 218.6639, 218.6632, 218.668, 218.6887, 218.6727, 218.6898, 218.6729, 218.6807, 218.6857, 218.6866, 218.6953, 218.6724, 218.6911, 218.6948, 218.6792, 218.68, 218.6922, 218.692, 218.6904, 218.6977, 218.7054, 218.6931, 218.7103, 218.6892, 218.6973, 218.6913, 218.6985, 218.7075, 218.6888, 218.6898, 218.6962, 218.6911, 218.6944, 218.7048, 218.7259, 218.7074, 218.6955, 218.6998, 218.7175, 218.699, 218.7068, 218.7252, 218.7222, 218.7167, 218.7361, 218.706, 218.7185, 218.7274, 218.7049, 218.7202, 218.7208, 218.7297, 218.748, 218.7209, 218.734, 218.7131, 218.7352, 218.7266, 218.7352, 218.7319, 218.7249, 218.7477, 218.7318, 218.7239, 218.7384, 218.7612, 218.7652, 218.7461, 218.7392, 218.7613, 218.75, 218.7701, 218.7572, 218.7641, 218.768, 218.7547, 218.7387, 218.7474, 218.7475, 218.754, 218.7769, 218.7707, 218.7596, 218.77, 218.7683, 218.7671, 218.7573, 218.7742, 218.7811, 218.7698, 218.7685, 218.7705, 218.7722, 218.7852, 218.7912, 218.798, 218.7791, 218.7969, 218.7892, 218.7699, 218.7856, 218.7733, 218.7953, 218.7939, 218.7935, 218.8021, 218.7982, 218.7776, 218.7873, 218.8031, 218.8016, 218.8089, 218.804, 218.791, 218.7918, 218.7947, 218.8061, 218.7955, 218.7997, 218.8003, 218.7963, 218.7896, 218.7912, 218.7897, 218.8097, 218.8122, 218.7991, 218.7914, 218.8111, 218.8049, 218.8113, 218.816, 218.8051, 218.8094, 218.813, 218.808, 218.8057, 218.808, 218.8169, 218.8087, 218.8085, 218.8173, 218.8191, 218.8082, 218.8197, 218.8093, 218.8099, 218.8169, 218.8132, 218.8169, 218.8024, 218.8351, 218.8164, 218.8033, 218.8191, 218.8081, 218.8181, 218.8161, 218.8103, 218.7959, 218.8251, 218.8004, 218.8298, 218.823, 218.8068, 218.8033, 218.8198, 218.7935, 218.8229, 218.8009, 218.8061, 218.815, 218.7956, 218.7972, 218.7914, 218.7905, 218.8023, 218.8009, 218.7991, 218.8123, 218.811, 218.8, 218.8061, 218.8026, 218.7955, 218.803, 218.8113, 218.7968, 218.8012, 218.8053, 218.8122, 218.7955, 218.7957, 218.7943, 218.7917, 218.7979, 218.7849, 218.8022, 218.8075, 218.7878, 218.7811, 218.783, 218.7926, 218.7915, 218.7817, 218.7907, 218.7856, 218.807, 218.7854, 218.8023, 218.8066, 218.8081, 218.7635, 218.7797, 218.7771, 218.7897, 218.7881, 218.7903, 218.7679, 218.7562, 218.7895, 218.766, 218.7598, 218.7606, 218.7632, 218.7585, 218.7813, 218.7637, 218.7441, 218.7487, 218.7657, 218.7497, 218.7531, 218.7607, 218.7417, 218.7599, 218.7513, 218.7504, 218.7387, 218.7334, 218.765, 218.7296, 218.7308, 218.7386, 218.7273, 218.7353, 218.735, 218.7354, 218.7258, 218.7107, 218.7354, 218.7112, 218.7049, 218.6943, 218.7071, 218.7093, 218.7002, 218.7002, 218.6754, 218.6899, 218.6778, 218.6871, 218.6778, 218.6752, 218.6852, 218.6833, 218.6743, 218.6665, 218.6727, 218.6802, 218.6699, 218.6623, 218.6688, 218.6708, 218.6608, 218.6501, 218.6508, 218.6463, 218.6517, 218.6404, 218.6476, 218.6356, 218.6418, 218.6388, 218.6363, 218.6251, 218.6362, 218.6163, 218.6275, 218.618, 218.6321, 218.6196, 218.6227, 218.6054, 218.5973, 218.6113, 218.5885, 218.6053, 218.6026, 218.5914, 218.5993, 218.5881, 218.5936, 218.592, 218.5911, 218.601, 218.6011, 218.585, 218.5701, 218.5822, 218.5739, 218.5722, 218.5789, 218.5671, 218.5687, 218.5546, 218.5649, 218.5639, 218.5566, 218.5477, 218.5504, 218.5361, 218.5412, 218.5228, 218.5349, 218.5493, 218.5499, 218.5298, 218.5263, 218.5369, 218.5307, 218.5237, 218.5167, 218.5279, 218.5225, 218.5171, 218.5129, 218.5154, 218.5133, 218.5146, 218.5203, 218.5011, 218.5102, 218.5142, 218.5006, 218.4804, 218.4905, 218.4914, 218.4966, 218.5056, 218.4785, 218.4915, 218.4624, 218.4722, 218.4816, 218.4891, 218.4704, 218.4827, 218.4547, 218.4722, 218.4736, 218.4712, 218.4523, 218.4748, 218.4502, 218.4546, 218.4597, 218.457, 218.4459, 218.4624, 218.4316, 218.4662, 218.4616, 218.4384, 218.4567, 218.4474, 218.4516, 218.448, 218.4343, 218.4475, 218.4565, 218.4483, 218.4358, 218.4192, 218.4463, 218.4402, 218.4446, 218.4193, 218.4303, 218.4339, 218.4288, 218.4269, 218.417, 218.4292, 218.4289, 218.4168, 218.4193, 218.4275, 218.4049, 218.411, 218.4189, 218.4076, 218.3958, 218.4066, 218.4137, 218.4049, 218.3993, 218.4034, 218.3917, 218.388, 218.4002, 218.3812, 218.4035, 218.3906, 218.3768, 218.4099, 218.4015, 218.3871, 218.3863, 218.3917, 218.3895, 218.3912, 218.3956, 218.3859, 218.3696, 218.3891, 218.3762, 218.3912, 218.3886, 218.3801, 218.3752, 218.39, 218.3656, 218.3884, 218.3806, 218.3771, 218.3881, 218.365, 218.3617, 218.388, 218.3653, 218.3864, 218.3727, 218.3743, 218.3838, 218.3722, 218.3732, 218.3718, 218.3799, 218.3893, 218.3971, 218.3896, 218.3826, 218.3845, 218.3858, 218.3883, 218.3934, 218.3873, 218.3867, 218.3877, 218.3975, 218.4016, 218.4099, 218.4061, 218.4344, 218.4151, 218.4323, 218.411, 218.4229, 218.4178, 218.4124, 218.4162, 218.4317, 218.4185, 218.4268, 218.417, 218.4194, 218.4374, 218.4384, 218.4378, 218.446, 218.4491, 218.4437, 218.4384, 218.4367, 218.4287, 218.4459, 218.4239, 218.438, 218.4463, 218.4461, 218.4544, 218.4495, 218.4547, 218.4354, 218.4428, 218.4513, 218.4562, 218.4464, 218.4473, 218.4432, 218.4521, 218.4443, 218.4584, 218.4496, 218.4516, 218.4575, 218.4476, 218.4426, 218.4456, 218.4465, 218.4575, 218.4607, 218.4639, 218.4634, 218.4609, 218.4482, 218.4658, 218.4672, 218.4505, 218.4498, 218.4495, 218.4666, 218.4616, 218.4703, 218.4598, 218.4745, 218.4652, 218.453, 218.4695, 218.4713, 218.454, 218.4736, 218.4694, 218.4706, 218.4752, 218.472, 218.4836, 218.4651, 218.4741, 218.4783, 218.4783, 218.4773, 218.4819, 218.4773, 218.4904, 218.4889, 218.4834, 218.4818, 218.4995, 218.4811, 218.4756, 218.478, 218.4811, 218.4913, 218.496, 218.4819, 218.4959, 218.5031, 218.5007, 218.496, 218.4932, 218.5007, 218.504, 218.4966, 218.4985, 218.5023, 218.5126, 218.5087, 218.5169, 218.5108, 218.5145, 218.5259, 218.5196, 218.5179, 218.5196, 218.526, 218.5105, 218.5198, 218.5204, 218.5082, 218.5236, 218.5202, 218.5264, 218.5223, 218.535, 218.5381, 218.5233, 218.5265, 218.5354, 218.5338, 218.5331, 218.5444, 218.5444, 218.5332, 218.5398, 218.5336, 218.5412, 218.5429, 218.5525, 218.5491, 218.5577, 218.5477, 218.5492, 218.5527, 218.5639, 218.5659, 218.5573, 218.5625, 218.563, 218.5535, 218.5602, 218.5659, 218.5527, 218.5763, 218.5688, 218.5592, 218.575, 218.5523, 218.5711, 218.5658, 218.5637, 218.5916, 218.579, 218.5639, 218.5841, 218.5772, 218.5859, 218.5897, 218.5914, 218.5871, 218.5851, 218.5949, 218.5889, 218.578, 218.592, 218.5961, 218.5949, 218.5953, 218.5835, 218.5952, 218.601, 218.6041, 218.6179, 218.5983, 218.6015, 218.6008, 218.6045, 218.6018, 218.6196, 218.6086, 218.6113, 218.6066, 218.6101, 218.6091, 218.6111, 218.6223, 218.6125, 218.6203, 218.6162, 218.6203, 218.6269, 218.6241, 218.6167, 218.6205, 218.6335, 218.6281, 218.6146, 218.6234, 218.6269, 218.6285, 218.6203, 218.6252, 218.6114, 218.6066, 218.6209, 218.6064, 218.6039, 218.5996, 218.5911, 218.6067, 218.6127, 218.6204, 218.6049, 218.6161, 218.6168, 218.6161, 218.621, 218.6105, 218.6231, 218.6203, 218.6286, 218.6266, 218.639, 218.6158, 218.6143, 218.6219, 218.633, 218.617, 218.6321, 218.6308, 218.6117, 218.6161, 218.6208, 218.6287, 218.6346, 218.6448, 218.6369, 218.6279, 218.6297, 218.6152, 218.625, 218.6418, 218.6283, 218.6254, 218.6428, 218.6407, 218.6203, 218.6255, 218.6241, 218.6346, 218.6362, 218.6395, 218.6374, 218.6534, 218.6779, 218.6793, 218.6736, 218.6778, 218.6888, 218.6801, 218.6875, 218.6918, 218.6866, 218.6959, 218.7028, 218.6866, 218.7025, 218.6941, 218.6959, 218.6908, 218.6898, 218.6877, 218.6844, 218.7073, 218.7026, 218.7215, 218.7037, 218.7116, 218.7096, 218.716, 218.7219, 218.715, 218.7274, 218.7317, 218.7234, 218.7242, 218.7164, 218.7105, 218.727, 218.7274, 218.7229, 218.7169, 218.7186, 218.7314, 218.7227, 218.7167, 218.7225, 218.7215, 218.7146, 218.73, 218.7209, 218.7296, 218.7471, 218.7379, 218.7522, 218.7377, 218.7544, 218.7607, 218.7464, 218.7569, 218.7486, 218.7614, 218.7656, 218.7732, 218.7657, 218.7652, 218.7685, 218.7768, 218.7808, 218.7749, 218.7744, 218.7745, 218.7744, 218.7761, 218.7954, 218.7839, 218.7881, 218.7852, 218.797, 218.7964, 218.7912, 218.7908, 218.8117, 218.8, 218.8048, 218.809, 218.8008, 218.8021, 218.8082, 218.8026, 218.8228, 218.8242, 218.8181, 218.8215, 218.8176, 218.8181, 218.8092, 218.8257, 218.8207, 218.831, 218.8251, 218.8264, 218.8178, 218.8291, 218.8223, 218.8295, 218.8316, 218.8446, 218.8257, 218.8411, 218.8552, 218.8285, 218.8586, 218.8469, 218.8504, 218.8447, 218.8628, 218.856, 218.8697, 218.8659, 218.8728, 218.8537, 218.8459, 218.8719, 218.8717, 218.848, 218.8739, 218.8691, 218.8712, 218.8697, 218.875, 218.8792, 218.8626, 218.8864, 218.8773, 218.88, 218.8821, 218.8832, 218.8785, 218.8967, 218.8931, 218.8818, 218.8765, 218.8933, 218.8886, 218.882, 218.8881, 218.8942, 218.8848, 218.8991, 218.8928, 218.8961, 218.8956, 218.8901, 218.8927, 218.8926, 218.8906, 218.8905, 218.8966, 218.902, 218.9027, 218.8862, 218.8846, 218.9061, 218.9043, 218.9021, 218.896, 218.9009, 218.8996, 218.9108, 218.902, 218.9027, 218.9014, 218.9132, 218.9061, 218.9152, 218.8989, 218.9037, 218.9181, 218.9058, 218.9119, 218.8906, 218.9147, 218.9265, 218.9229, 218.9021, 218.9189, 218.9151, 218.9057, 218.9125, 218.8977, 218.9007, 218.9167, 218.9101, 218.9031, 218.9101, 218.9081, 218.9177, 218.9086, 218.9133, 218.9133, 218.9097, 218.914, 218.8984, 218.908, 218.9078, 218.8979, 218.9081, 218.9093, 218.8982, 218.9075, 218.8982, 218.8837, 218.8841, 218.8897, 218.8934, 218.8867, 218.888, 218.8863, 218.8831, 218.883, 218.8747, 218.8832, 218.8866, 218.8728, 218.886, 218.8703, 218.864, 218.8614, 218.8557, 218.8755, 218.8646, 218.833, 218.8514, 218.8441, 218.8586, 218.8508, 218.8549, 218.8366, 218.8357, 218.8347, 218.8402, 218.822, 218.8403, 218.8123, 218.8102, 218.8105, 218.804, 218.8121, 218.7973, 218.7906, 218.8102, 218.7936, 218.8008, 218.8022, 218.7978, 218.7855, 218.7694, 218.7903, 218.7922, 218.7714, 218.7668, 218.7897, 218.7845, 218.775, 218.7584, 218.7713, 218.7748, 218.7638, 218.7527, 218.7702, 218.7641, 218.7594, 218.7531, 218.7445, 218.7504, 218.7335, 218.7433, 218.734, 218.7164, 218.7275, 218.7059, 218.7114, 218.6966, 218.6912, 218.7063, 218.6927, 218.6915, 218.6957, 218.6941, 218.6828, 218.6846, 218.6965, 218.6755, 218.6692, 218.6692, 218.653, 218.6638, 218.6807, 218.6604, 218.6555, 218.6587, 218.6511, 218.6342, 218.6463, 218.6413, 218.6194, 218.6365, 218.6328, 218.6286, 218.6348, 218.6105, 218.6126, 218.609, 218.609, 218.6129, 218.6163, 218.6087, 218.6149, 218.5903, 218.5773, 218.5927, 218.5992, 218.588, 218.5788, 218.583, 218.5824, 218.5702, 218.5601, 218.5643, 218.5692, 218.5688, 218.5455, 218.5587, 218.5562, 218.5519, 218.5522, 218.5462, 218.5545, 218.5367, 218.5344, 218.5254, 218.5337, 218.5159, 218.5218, 218.5172, 218.5121, 218.5073, 218.509, 218.5083, 218.51, 218.5155, 218.5029, 218.5095, 218.4925, 218.5063, 218.4901, 218.4842, 218.4663, 218.4968, 218.4829, 218.4899, 218.4858, 218.4826, 218.4775, 218.4738, 218.4512, 218.4863, 218.4743, 218.4534, 218.461, 218.4658, 218.4619, 218.4608, 218.4524, 218.4539, 218.4459, 218.4477, 218.4512, 218.4448, 218.4488, 218.4467, 218.4451, 218.4448, 218.4482, 218.4275, 218.4403, 218.4359, 218.4433, 218.4272, 218.4298, 218.4341, 218.4295, 218.4196, 218.4124, 218.4206, 218.4162, 218.4192, 218.4175, 218.4135, 218.4041, 218.4102, 218.4276, 218.4074, 218.4122, 218.4054, 218.4094, 218.3914, 218.3922, 218.4036, 218.3898, 218.3994, 218.4032, 218.3865, 218.3782, 218.4, 218.3953, 218.3711, 218.3849, 218.3774, 218.393, 218.3901, 218.3877, 218.3831, 218.3618, 218.3737, 218.3827, 218.388, 218.3698, 218.3724, 218.3664, 218.3817, 218.3724, 218.3595, 218.3745, 218.3682, 218.3577, 218.3662, 218.3541, 218.367, 218.3707, 218.368, 218.3714, 218.3753, 218.3655, 218.3689, 218.3657, 218.367, 218.3598, 218.3729, 218.3688, 218.3739, 218.3726, 218.3578, 218.3753, 218.3669, 218.3654, 218.3899, 218.3563, 218.3697, 218.3729, 218.3735, 218.3654, 218.3638, 218.3638, 218.3842, 218.3769, 218.377, 218.3826, 218.3732, 218.3821, 218.3754, 218.3669, 218.3743, 218.3771, 218.3933, 218.3776, 218.3943, 218.3868, 218.3981, 218.4, 218.3849, 218.396, 218.3877, 218.3918, 218.3848, 218.3956, 218.3842, 218.4043, 218.3868, 218.3933, 218.4018, 218.4022, 218.384, 218.3791, 218.3986, 218.4114, 218.4022, 218.4065, 218.4065, 218.4011, 218.4004, 218.4156, 218.4035, 218.4082, 218.4019, 218.4126, 218.4128, 218.4165, 218.4191, 218.41, 218.4104, 218.4035, 218.4345, 218.4207, 218.4176, 218.4252, 218.4137, 218.4214, 218.425, 218.418, 218.4282, 218.4213, 218.4251, 218.4399, 218.4146, 218.4178, 218.4263, 218.4173, 218.4496, 218.4338, 218.4204, 218.4408, 218.4345, 218.448, 218.438, 218.4327, 218.4344, 218.4488, 218.448, 218.4555, 218.4398, 218.4551, 218.4613, 218.4581, 218.4553, 218.4659, 218.4689, 218.4594, 218.4725, 218.4642, 218.4584, 218.4583, 218.48, 218.4685, 218.4774, 218.4635, 218.4693, 218.4757, 218.476, 218.4691, 218.4805, 218.4732, 218.4802, 218.4769, 218.4821, 218.4857, 218.4689, 218.4882, 218.4909, 218.4791, 218.4819, 218.4889, 218.5006, 218.5028, 218.5022, 218.488, 218.4969, 218.5037, 218.4933, 218.4971, 218.4995, 218.5009, 218.5084, 218.518, 218.5106, 218.5199, 218.514, 218.5373, 218.521, 218.5232, 218.52, 218.5433, 218.5335, 218.5301, 218.5325, 218.5347, 218.5413, 218.5304, 218.5455, 218.5394, 218.5466, 218.5289, 218.5437, 218.5505, 218.552, 218.5457, 218.5593, 218.5533, 218.5651, 218.5652, 218.5505, 218.5593, 218.5607, 218.5788, 218.5734, 218.5732, 218.5712, 218.5824, 218.5727, 218.5841, 218.5737, 218.576, 218.5873, 218.586, 218.5806, 218.5881, 218.5853, 218.5866, 218.5888, 218.5922, 218.5988, 218.606, 218.5914, 218.5857, 218.6004, 218.608, 218.5949, 218.5993, 218.6032, 218.6076, 218.5995, 218.6071, 218.6077, 218.6213, 218.613, 218.6062, 218.6129, 218.6003, 218.6081, 218.614, 218.6137, 218.6139, 218.6139, 218.6244, 218.613, 218.6017, 218.6184, 218.6091, 218.6137, 218.6197, 218.6045, 218.6105, 218.6139, 218.6324, 218.6228, 218.6234, 218.6338, 218.626, 218.6263, 218.639, 218.6344, 218.6489, 218.6318, 218.6469, 218.6338, 218.6465, 218.637, 218.6526, 218.6528, 218.6376, 218.6514, 218.644, 218.6571, 218.6355, 218.6385, 218.6304, 218.6483, 218.6528, 218.6534, 218.6493, 218.6419, 218.6598, 218.6484, 218.6639, 218.6618, 218.6759, 218.6722, 218.6576, 218.6658, 218.6593, 218.6531, 218.659, 218.6693, 218.6749, 218.6614, 218.6662, 218.6731, 218.6693, 218.6681, 218.6712, 218.6655, 218.6807, 218.6792, 218.6729, 218.675, 218.6847, 218.6789, 218.6939, 218.6934, 218.6751, 218.6764, 218.6801, 218.6861, 218.6962, 218.7008, 218.6954, 218.7091, 218.7082, 218.6834, 218.7009, 218.6969, 218.6944, 218.6928, 218.6945, 218.6818, 218.7093, 218.7, 218.7135, 218.7032, 218.711, 218.7256, 218.7092, 218.7281, 218.7107, 218.7212, 218.7256, 218.7086, 218.7252, 218.7154, 218.7236, 218.734, 218.7155, 218.7477, 218.7302, 218.7206, 218.7303, 218.7333, 218.7339, 218.7425, 218.7443, 218.7537, 218.734, 218.7481, 218.7474, 218.754, 218.7536, 218.7713, 218.7703, 218.7625, 218.7648, 218.778, 218.7806, 218.7719, 218.7724, 218.7735, 218.7852, 218.7997, 218.7874, 218.7894, 218.8006, 218.7852, 218.8059, 218.81, 218.817, 218.8071, 218.809, 218.8038, 218.8122, 218.8133, 218.8018, 218.8116, 218.8028, 218.8201, 218.8195, 218.8356, 218.8335, 218.8255, 218.8257, 218.8289, 218.8245, 218.8261, 218.8292, 218.8297, 218.836, 218.8401, 218.8395, 218.844, 218.8477, 218.8504, 218.8562, 218.8682, 218.8666, 218.8585, 218.8633, 218.8467, 218.8734, 218.8594, 218.8813, 218.8627, 218.8723, 218.8792, 218.8854, 218.8851, 218.8685, 218.8779, 218.8764, 218.8936, 218.8765, 218.8841, 218.8827, 218.8851, 218.883, 218.8933, 218.8946, 218.9029, 218.8974, 218.9078, 218.9147, 218.9133, 218.9125, 218.9086, 218.908, 218.9206, 218.9356, 218.9315, 218.9252, 218.9172, 218.9325, 218.9243, 218.9394, 218.9262, 218.9288, 218.9407, 218.9374, 218.9514, 218.9433, 218.9445, 218.9472, 218.9567, 218.942, 218.9653, 218.9549, 218.9541, 218.9557, 218.9558, 218.9722, 218.9677, 218.9592, 218.9626, 218.9769, 218.9777, 218.9853, 218.9751, 218.9825, 218.9831, 218.9862, 218.9849, 218.993, 219.0037, 218.9892, 218.9948, 218.9909, 218.9916, 218.9801, 218.9973, 218.9848, 218.9959, 218.9836, 219.0077, 219.0067, 218.9916, 218.9894, 219.0118, 219.0102, 219.0035, 219.0112, 219.0086, 218.9964, 219.0011, 219.0052, 219.0035, 219.0126, 219.0071, 219.0206, 219.0159, 219.0189, 219.0224, 219.0124, 219.0137, 219.0133, 219.0086, 219.0027, 219.0192, 219.0078, 219.0153, 218.9979, 219.007, 218.9953, 219.0049, 218.9879, 219.0238, 219.0088, 219.0032, 219.0255, 219.0067, 219.0095, 218.9907, 218.9943, 218.9978, 218.9969, 219.0105, 218.9859, 218.9908, 219.0055, 218.9978, 218.969, 219.0026, 218.9939, 218.9944, 218.9831, 218.9759, 218.9777, 218.9859, 218.9644, 218.9819, 218.972, 218.9515, 218.9595, 218.9567, 218.952, 218.9615, 218.9511, 218.9593, 218.942, 218.9529, 218.9441, 218.9435, 218.9419, 218.9415, 218.9335, 218.9308, 218.9285, 218.9447, 218.93, 218.9282, 218.9442, 218.92, 218.9213, 218.9166, 218.9261, 218.9323, 218.9226, 218.8963, 218.9232, 218.9145, 218.9089, 218.9026, 218.8788, 218.8848, 218.897, 218.8869, 218.8877, 218.8739, 218.8725, 218.8656, 218.8657, 218.8775, 218.8553, 218.877, 218.8562, 218.8563, 218.8506, 218.8498, 218.8445, 218.8393, 218.8256, 218.8258, 218.8238, 218.8306, 218.8177, 218.8197, 218.8231, 218.8077, 218.8171, 218.8135, 218.8015, 218.804, 218.7995, 218.7955, 218.7929, 218.7835, 218.7939, 218.7855, 218.7633, 218.7652, 218.7693, 218.7647, 218.759, 218.7568, 218.7563, 218.7456, 218.7634, 218.7487, 218.7372, 218.7375, 218.7396, 218.7307, 218.7233, 218.7114, 218.7089, 218.71, 218.7001, 218.696, 218.7042, 218.6852, 218.698, 218.6921, 218.6777, 218.6866, 218.6586, 218.6607, 218.6652, 218.6652, 218.6644, 218.6535, 218.6482, 218.6432, 218.6528, 218.6513, 218.6212, 218.636, 218.6392, 218.6277, 218.6205, 218.6068, 218.6199, 218.6107, 218.6169, 218.6067, 218.6067, 218.6041, 218.6005, 218.5857, 218.5922, 218.5956, 218.5876, 218.5768, 218.5872, 218.5769, 218.5648, 218.5586, 218.5639, 218.5693, 218.5488, 218.5629, 218.5463, 218.5744, 218.5511, 218.5466, 218.5509, 218.5509, 218.532, 218.5222, 218.5257, 218.5345, 218.5279, 218.5114, 218.5118, 218.5171, 218.5044, 218.4846, 218.4887, 218.4965, 218.4884, 218.4675, 218.4976, 218.497, 218.4839, 218.5098, 218.4917, 218.4687, 218.4715, 218.4684, 218.4615, 218.4719, 218.4581, 218.4645, 218.4405, 218.463, 218.4526, 218.4461, 218.4427, 218.4301, 218.4371, 218.4259, 218.4467, 218.4253, 218.4207, 218.4339, 218.4433, 218.4433, 218.4108, 218.4124, 218.4276, 218.3937, 218.4245, 218.4023, 218.3933, 218.3965, 218.3958, 218.4069, 218.4191, 218.4017, 218.421, 218.41, 218.3843, 218.4012, 218.3937, 218.3906, 218.3835, 218.3855, 218.3827, 218.3912, 218.3772, 218.3661, 218.3807, 218.3798, 218.3874, 218.3716, 218.3826, 218.362, 218.3645, 218.3669, 218.3658, 218.3486, 218.3565, 218.375, 218.3835, 218.376, 218.354, 218.3463, 218.3511, 218.3661, 218.3364, 218.3544, 218.3462, 218.3496, 218.3548, 218.3306, 218.3741, 218.3466, 218.3457, 218.3555, 218.3457, 218.3418, 218.3414, 218.3561, 218.3385, 218.3327, 218.3258, 218.3413, 218.3393, 218.3474, 218.3403, 218.3414, 218.334, 218.3453, 218.333, 218.3289, 218.3375, 218.3337, 218.3384, 218.3352, 218.3434, 218.346, 218.3413, 218.3416, 218.3624, 218.3304, 218.3365, 218.3596, 218.3475, 218.355, 218.3669, 218.3686, 218.3499, 218.3453, 218.3469, 218.3499, 218.3631, 218.3825, 218.3607, 218.3555, 218.3749, 218.3711, 218.3667, 218.3512, 218.3635, 218.3757, 218.3784, 218.3709, 218.374, 218.3684, 218.3714, 218.3679, 218.3772, 218.3831, 218.3909, 218.3856, 218.3889, 218.3795, 218.3947, 218.3873, 218.3953, 218.3885, 218.394, 218.4191, 218.3971, 218.4056, 218.3906, 218.4054, 218.4059, 218.3987, 218.4213, 218.3959, 218.4042, 218.424, 218.4343, 218.4112, 218.4176, 218.4229, 218.4111, 218.422, 218.4308, 218.43, 218.4347, 218.4344, 218.4197, 218.42, 218.4464, 218.4206, 218.4427, 218.4401, 218.4319, 218.4335, 218.4406, 218.4405, 218.4474, 218.454, 218.4436, 218.4646, 218.4558, 218.4588, 218.4644, 218.4614, 218.4333, 218.4838, 218.4644, 218.4596, 218.4842, 218.4886, 218.4948, 218.4773, 218.514, 218.4959, 218.4787, 218.4832, 218.4937, 218.4874, 218.4956, 218.5166, 218.498, 218.5064, 218.5178, 218.5061, 218.5186, 218.504, 218.5148, 218.5202, 218.5062, 218.4944, 218.5179, 218.5338, 218.52, 218.5309, 218.537, 218.5331, 218.51, 218.5337, 218.5352, 218.5147, 218.5606, 218.5483, 218.5374, 218.5467, 218.561, 218.5693, 218.5637, 218.5482, 218.5543, 218.5644, 218.5611, 218.5667, 218.5383, 218.5477, 218.5562, 218.5592, 218.5704, 218.5427, 218.5847, 218.5621, 218.5556, 218.5744, 218.5794, 218.5798, 218.5936, 218.5894, 218.5699, 218.5704, 218.5832, 218.5782, 218.6082, 218.5889, 218.5879, 218.5928, 218.5927, 218.5912, 218.618, 218.613, 218.615, 218.5989, 218.5869, 218.5846, 218.6158, 218.6046, 218.5903, 218.6216, 218.6144, 218.5815, 218.5907, 218.6039, 218.6074, 218.614, 218.6008, 218.5994, 218.62, 218.6319, 218.6285, 218.617, 218.6212, 218.6205, 218.6463, 218.6148, 218.6118, 218.606, 218.6258, 218.6457, 218.6605, 218.6522, 218.6479, 218.6347, 218.6284, 218.6374, 218.6402, 218.6381, 218.6567, 218.6511, 218.6331, 218.6403, 218.627, 218.6098, 218.6102, 218.6224, 218.6322, 218.6416, 218.6322, 218.6424, 218.6434, 218.6365, 218.6694, 218.666, 218.6272, 218.6523, 218.6609, 218.6633, 218.6705, 218.6829, 218.6534, 218.6644, 218.657, 218.678, 218.6623, 218.6593, 218.6421, 218.6667, 218.6676, 218.6563, 218.6647, 218.6571, 218.6653, 218.6847, 218.6675, 218.6871, 218.6765, 218.6931, 218.6745, 218.6797, 218.6735, 218.6803, 218.6693, 218.6795, 218.6664, 218.6746, 218.6896, 218.6815, 218.6851, 218.6721, 218.7017, 218.6874, 218.695, 218.7019, 218.6795, 218.6983, 218.7121, 218.6998, 218.6922, 218.7061, 218.689, 218.6865, 218.6863, 218.6844, 218.6891, 218.7091, 218.7021, 218.6969, 218.6953, 218.7022, 218.6953, 218.6782, 218.7126, 218.6976, 218.6877, 218.7276, 218.7, 218.7004, 218.7215, 218.727, 218.6916, 218.7024, 218.7163, 218.7412, 218.7142, 218.7235, 218.7157, 218.7036, 218.71, 218.7188, 218.7282, 218.7269, 218.7176, 218.7283, 218.7386, 218.7513, 218.7269, 218.7317, 218.7268, 218.7544, 218.7235, 218.7243, 218.7356, 218.739, 218.7381, 218.7693, 218.7623, 218.7542, 218.7484, 218.7605, 218.7689, 218.7701, 218.7818, 218.7799, 218.7875, 218.7919, 218.7766, 218.7978, 218.7829, 218.7769, 218.7895, 218.7923, 218.7997, 218.8046, 218.8103, 218.7998, 218.806, 218.8154, 218.8235, 218.8256, 218.82, 218.8308, 218.8288, 218.815, 218.8214, 218.8496, 218.8346, 218.8279, 218.8327, 218.8434, 218.8369, 218.8436, 218.8637, 218.8423, 218.8422, 218.8416, 218.851, 218.8592, 218.8696, 218.8725, 218.8813, 218.8868, 218.8563, 218.8622, 218.886, 218.8831, 218.8717, 218.88, 218.8866, 218.8961, 218.8846, 218.9034, 218.903, 218.8974, 218.9008, 218.9118, 218.9085, 218.9193, 218.9194, 218.9188, 218.9062, 218.9384, 218.9241, 218.913, 218.9347, 218.9394, 218.9207, 218.9275, 218.9306, 218.9326, 218.9331, 218.9514, 218.9397, 218.944, 218.9366, 218.9454, 218.9557, 218.9643, 218.9534, 218.9667, 218.9615, 218.9617, 218.9673, 218.9756, 218.9772, 218.9874, 218.9766, 218.9795, 218.9937, 218.9906, 218.9752, 218.9888, 218.9813, 218.9999, 218.9726, 218.9995, 219.0001, 218.9967, 218.9978, 219.0109, 219.0116, 219.013, 219.0106, 219.0168, 219.0064, 219.0222, 218.9987, 219.0419, 219.0212, 219.0288, 219.0208, 219.0315, 219.0309, 219.022, 219.0337, 219.0259, 219.0284, 219.0482, 219.0355, 219.0189, 219.0273, 219.044, 219.0536, 219.0425, 219.0477, 219.0589, 219.0547, 219.0444, 219.06, 219.043, 219.057, 219.0448, 219.0475, 219.0566, 219.0678, 219.0516, 219.0537, 219.0443, 219.0677, 219.0523, 219.0536, 219.0574, 219.0713, 219.0815, 219.0661, 219.065, 219.0764, 219.0502, 219.0882, 219.0548, 219.0675, 219.0841, 219.0541, 219.0805, 219.0779, 219.0577, 219.0619, 219.0592, 219.061, 219.0777, 219.0583, 219.0798, 219.0614, 219.0723, 219.0635, 219.0784, 219.0627, 219.0722, 219.0609, 219.0514, 219.0621, 219.0526, 219.0736, 219.0668, 219.0558, 219.0562, 219.0546, 219.0588, 219.024, 219.0411, 219.0467, 219.0478, 219.048, 219.0214, 219.0364, 219.0189, 219.0421, 219.0215, 219.036, 219.0267, 219.0192, 219.0186, 219.0137, 219.0171, 219.0277, 219.0023, 218.9956, 218.9962, 219.0224, 218.9833, 218.9852, 218.996, 218.9804, 218.9917, 218.9963, 218.9943, 218.9948, 218.9722, 218.9783, 218.9708, 218.975, 218.9661, 218.952, 218.9598, 218.9678, 218.9385, 218.9425, 218.948, 218.9571, 218.9305, 218.95, 218.9285, 218.915, 218.9156, 218.924, 218.919, 218.9023, 218.9181, 218.903, 218.9259, 218.9048, 218.8966, 218.8814, 218.8962, 218.8694, 218.903, 218.884, 218.8658, 218.8993, 218.8732, 218.8698, 218.8569, 218.8553, 218.8435, 218.8442, 218.8467, 218.8591, 218.8499, 218.8411, 218.8424, 218.8258, 218.8285, 218.831, 218.7872, 218.8273, 218.794, 218.8098, 218.7877, 218.7961, 218.8018, 218.7966, 218.7874, 218.7839, 218.7834, 218.7535, 218.7789, 218.7645, 218.7603, 218.7588, 218.755, 218.7516, 218.7471, 218.739, 218.7403, 218.7117, 218.7157, 218.7214, 218.7173, 218.7145, 218.7064, 218.7126, 218.7015, 218.6865, 218.7, 218.7055, 218.6864, 218.6712, 218.6908, 218.6811, 218.6434, 218.6859, 218.6689, 218.6592, 218.648, 218.6665, 218.6363, 218.6369, 218.661, 218.6412, 218.6403, 218.6337, 218.6186, 218.6229, 218.6293, 218.6202, 218.6179, 218.6136, 218.6032, 218.6025, 218.5962, 218.5881, 218.591, 218.6001, 218.5719, 218.5724, 218.5587, 218.5696, 218.5765, 218.551, 218.5558, 218.5586, 218.5643, 218.5446, 218.5436, 218.5329, 218.5219, 218.5452, 218.5154, 218.5349, 218.5341, 218.5202, 218.5313, 218.5127, 218.5149, 218.492, 218.5039, 218.4738, 218.5047, 218.5063, 218.4748, 218.4542, 218.4892, 218.4767, 218.4578, 218.4539, 218.4615, 218.4499, 218.4518, 218.4633, 218.4584, 218.4377, 218.4373, 218.4331, 218.4216, 218.4367, 218.4305, 218.4216, 218.4248, 218.4369, 218.4266, 218.4005, 218.4185, 218.3981, 218.4223, 218.4051, 218.4049, 218.4101, 218.3967, 218.379, 218.3968, 218.4022, 218.3797, 218.3789, 218.3999, 218.3826, 218.3884, 218.3672, 218.3876, 218.3799, 218.3742, 218.364, 218.365, 218.3651, 218.3663, 218.3655, 218.3553, 218.3714, 218.3952, 218.3646, 218.3519, 218.3626, 218.3719, 218.3708, 218.3422, 218.3563, 218.3573, 218.3541, 218.3797, 218.353, 218.3588, 218.3737, 218.3472, 218.3447, 218.3701, 218.375, 218.3694, 218.3456, 218.3592, 218.3634, 218.3587, 218.3655, 218.3452, 218.3525, 218.3452, 218.3651, 218.3644, 218.3548, 218.3577, 218.3551, 218.3362, 218.3678, 218.3468, 218.3517, 218.3518, 218.3556, 218.3607, 218.3452, 218.3311, 218.3528, 218.3455, 218.3489, 218.3486, 218.3524, 218.3587, 218.3677, 218.3609, 218.3619, 218.3501, 218.3356, 218.3656, 218.3416, 218.3358, 218.3543, 218.3475, 218.3606, 218.3537, 218.3575, 218.3496, 218.358, 218.3666, 218.3463, 218.3701, 218.3635, 218.3701, 218.3664, 218.3672, 218.3711, 218.3603, 218.3774, 218.3776, 218.3803, 218.3855, 218.3831, 218.3691, 218.3736, 218.3876, 218.3799, 218.3975, 218.3774, 218.3864, 218.3867, 218.3792, 218.3905, 218.4046, 218.4024, 218.4052, 218.3976, 218.4026, 218.4045, 218.4167, 218.4027, 218.4118, 218.4264, 218.4158, 218.4159, 218.4213, 218.4128, 218.4277, 218.4241, 218.4065, 218.4272, 218.4314, 218.4221, 218.4317, 218.4203, 218.4298, 218.4358, 218.4444, 218.4473, 218.4426, 218.4455, 218.4474, 218.4568, 218.4367, 218.4429, 218.4461, 218.4332, 218.4682, 218.4376, 218.4489, 218.4379, 218.4694, 218.4665, 218.4762, 218.478, 218.476, 218.4834, 218.4788, 218.4886, 218.4671, 218.4914, 218.5084, 218.506, 218.5057, 218.514, 218.507, 218.5015, 218.4993, 218.5094, 218.5001, 218.5114, 218.5204, 218.5316, 218.5221, 218.5278, 218.5338, 218.5241, 218.5188, 218.5212, 218.5159, 218.5242, 218.5251, 218.5407, 218.553, 218.5286, 218.5524, 218.5471, 218.5438, 218.5493, 218.5456, 218.543, 218.5659, 218.5558, 218.5567, 218.5658, 218.5786, 218.5723, 218.5605, 218.5539, 218.5629, 218.5653, 218.5545, 218.5687, 218.5561, 218.5492, 218.5875, 218.568, 218.5724, 218.5787, 218.5788, 218.5728, 218.575, 218.5844, 218.5871, 218.5887, 218.585, 218.579, 218.6004, 218.596, 218.5895, 218.604, 218.5789, 218.5898, 218.6088, 218.6037, 218.6085, 218.6008, 218.5919, 218.5989, 218.6043, 218.6147, 218.6169, 218.6083, 218.6032, 218.6131, 218.6127, 218.6076, 218.5992, 218.6113, 218.5859, 218.603, 218.6018, 218.5977, 218.608, 218.624, 218.6221, 218.6155, 218.6292, 218.624, 218.6182, 218.6233, 218.6117, 218.6241, 218.6385, 218.6431, 218.6303, 218.6308, 218.6425, 218.6237, 218.624, 218.6323, 218.6252, 218.6413, 218.6338, 218.62, 218.6312, 218.6258, 218.6164, 218.6328, 218.6271, 218.641, 218.6331, 218.6303, 218.6152, 218.6231, 218.6269, 218.6353, 218.636, 218.6092, 218.6222, 218.6353, 218.6375, 218.6315, 218.6367, 218.6108, 218.6249, 218.625, 218.6013, 218.6253, 218.6274, 218.6318, 218.6443, 218.6405, 218.6412, 218.6388, 218.6419, 218.6153, 218.6227, 218.6353, 218.6296, 218.6472, 218.6382, 218.6454, 218.6388, 218.6406, 218.6414, 218.6442, 218.6418, 218.6485, 218.6345, 218.6548, 218.6584, 218.6338, 218.6304, 218.631, 218.6384, 218.6413, 218.6735, 218.6713, 218.6676, 218.6402, 218.6605, 218.6667, 218.6339, 218.6567, 218.6476, 218.647, 218.6536, 218.6674, 218.6762, 218.6896, 218.6734, 218.6724, 218.6693, 218.677, 218.6658, 218.6891, 218.6864, 218.6788, 218.6809, 218.6833, 218.6792, 218.7067, 218.7062, 218.6926, 218.6869, 218.7033, 218.6926, 218.7019, 218.7088, 218.7205, 218.7046, 218.7009, 218.7044, 218.7084, 218.717, 218.7089, 218.7065, 218.7154, 218.7305, 218.7388, 218.7292, 218.7099, 218.7418, 218.7292, 218.7277, 218.7278, 218.7407, 218.7313, 218.7446, 218.7477, 218.7462, 218.739, 218.7377, 218.7449, 218.7575, 218.7833, 218.7488, 218.7551, 218.7528, 218.7437, 218.7491, 218.7577, 218.7565, 218.7567, 218.7572, 218.7775, 218.7772, 218.7923, 218.7603, 218.7697, 218.7777, 218.8071, 218.7909, 218.7959, 218.8013, 218.809, 218.799, 218.7947, 218.8041, 218.8305, 218.8271, 218.82, 218.8187, 218.8291, 218.8446, 218.8264, 218.8369, 218.834, 218.8355, 218.8388, 218.8568, 218.8646, 218.8534, 218.8443, 218.8474, 218.8677, 218.8691, 218.863, 218.8773, 218.8804, 218.8913, 218.8752, 218.8835, 218.878, 218.8832, 218.9081, 218.891, 218.8975, 218.8994, 218.9022, 218.9031, 218.8998, 218.9137, 218.9015, 218.915, 218.9407, 218.9264, 218.9376, 218.9278, 218.9432, 218.9304, 218.9421, 218.9399, 218.9616, 218.9743, 218.9395, 218.9367, 218.9298, 218.9419, 218.9481, 218.9491, 218.9656, 218.9494, 218.945, 218.9614, 218.9596, 218.9754, 218.9613, 218.981, 218.9966, 219.0032, 218.9869, 218.9893, 218.9775, 218.9938, 218.9815, 218.9998, 219.008, 218.9954, 219.0029, 219.011, 219.0063, 219.0105, 218.9907, 219.0191, 219.0189, 219.0026, 219.0202, 219.0035, 219.0246, 219.0246, 219.0094, 219.0323, 219.0404, 219.0277, 219.0314, 219.0279, 219.0328, 219.0502, 219.0473, 219.0553, 219.0368, 219.0253, 219.0359, 219.0515, 219.0509, 219.0568, 219.0524, 219.0616, 219.0791, 219.0742, 219.0654, 219.0667, 219.0361, 219.0764, 219.0724, 219.078, 219.0488, 219.0685, 219.0547, 219.0701, 219.06, 219.0661, 219.0679, 219.091, 219.0814, 219.0455, 219.0649, 219.0877, 219.0713, 219.0712, 219.0911, 219.0732, 219.0722, 219.0742, 219.0724, 219.0742, 219.0796, 219.0673, 219.0622, 219.0648, 219.066, 219.066, 219.0625, 219.0789, 219.0655, 219.0771, 219.0673, 219.0908, 219.0582, 219.0689, 219.088, 219.076, 219.0657, 219.0762, 219.0837, 219.0669, 219.0578, 219.0532, 219.0614, 219.0472, 219.0558, 219.0774, 219.0668, 219.0482, 219.0318, 219.049, 219.0457, 219.0503, 219.0519, 219.035, 219.046, 219.0448, 219.0498, 219.0387, 219.0415, 219.0299, 219.0376, 219.0426, 219.0227, 219.0148, 219.0291, 219.0213, 219.0096, 219.0205, 219.0202, 219.0036, 219.021, 218.9945, 219.0125, 218.9996, 219.0103, 218.9981, 219.0146, 219.0165, 218.9929, 218.9962, 218.9841, 218.9846, 218.9893, 218.9802, 218.9544, 218.9848, 218.9569, 218.9848, 218.9595, 218.969, 218.9471, 218.9617, 218.9357, 218.9384, 218.9488, 218.9306, 218.908, 218.9252, 218.9308, 218.9223, 218.9098, 218.8985, 218.9139, 218.9076, 218.9104, 218.8924, 218.8996, 218.8891, 218.8985, 218.8802, 218.8672, 218.8646, 218.8927, 218.8748, 218.8422, 218.8696, 218.8483, 218.8597, 218.8549, 218.825, 218.8355, 218.8344, 218.8215, 218.817, 218.8274, 218.8109, 218.8052, 218.8078, 218.7968, 218.8138, 218.7925, 218.7678, 218.7827, 218.7819, 218.7756, 218.7725, 218.7763, 218.7663, 218.7652, 218.7281, 218.7519, 218.7383, 218.732, 218.7397, 218.7224, 218.725, 218.7161, 218.7075, 218.6929, 218.7053, 218.6896, 218.6805, 218.7141, 218.7105, 218.6749, 218.6765, 218.6686, 218.6708, 218.6529, 218.6535, 218.6605, 218.6607, 218.6702, 218.6418, 218.6407, 218.6333, 218.6023, 218.6333, 218.623, 218.5951, 218.6194, 218.6063, 218.6192, 218.5823, 218.5882, 218.6026, 218.5881, 218.5832, 218.5765, 218.5865, 218.5894, 218.5857, 218.563, 218.5723, 218.5724, 218.5448, 218.5511, 218.5352, 218.5354, 218.5219, 218.5508, 218.5345, 218.5352, 218.5036, 218.5257, 218.4908, 218.5231, 218.5023, 218.4995, 218.5073, 218.5152, 218.5125, 218.4736, 218.4966, 218.4737, 218.4763, 218.4731, 218.4748, 218.4501, 218.4683, 218.4547, 218.4782, 218.4523, 218.4647, 218.4533, 218.4659, 218.4436, 218.4473, 218.44, 218.4364, 218.4202, 218.4357, 218.432, 218.4117, 218.4305, 218.3836, 218.4056, 218.388, 218.412, 218.3936, 218.4013, 218.3766, 218.4004, 218.3986, 218.3866, 218.3792, 218.3872, 218.3859, 218.361, 218.3763, 218.3865, 218.3674, 218.3978, 218.3649, 218.3728, 218.3607, 218.3595, 218.3656, 218.3667, 218.3503, 218.3597, 218.366, 218.3557, 218.3493, 218.3455, 218.3382, 218.3674, 218.3563, 218.3477, 218.3478, 218.3551, 218.3715, 218.353, 218.3557, 218.3179, 218.3468, 218.338, 218.3438, 218.346, 218.33, 218.3342, 218.3559, 218.3217, 218.3352, 218.3215, 218.3264, 218.3153, 218.3366, 218.3386, 218.3191, 218.3142, 218.3236, 218.3141, 218.3262, 218.3018, 218.3105, 218.3289, 218.2998, 218.32, 218.3552, 218.3135, 218.3001, 218.314, 218.3307, 218.3002, 218.3095, 218.3122, 218.3298, 218.3468, 218.3289, 218.3183, 218.3364, 218.3432, 218.3288, 218.3372, 218.3262, 218.322, 218.3338, 218.327, 218.3405, 218.3141, 218.3297, 218.3283, 218.3183, 218.361, 218.3386, 218.3434, 218.3496, 218.3217, 218.3418, 218.3451, 218.3502, 218.3525, 218.333, 218.332, 218.3524, 218.3559, 218.3594, 218.365, 218.3625, 218.3642, 218.3773, 218.3631, 218.3652, 218.3566, 218.3713, 218.3766, 218.3922, 218.3809, 218.3725, 218.3572, 218.394, 218.3933, 218.414, 218.3875, 218.3798, 218.3945, 218.386, 218.3984, 218.3911, 218.387, 218.3965, 218.4157, 218.4197, 218.4027, 218.3784, 218.3918, 218.405, 218.416, 218.4092, 218.4153, 218.4103, 218.4137, 218.4198, 218.4362, 218.4198, 218.4198, 218.4128, 218.4301, 218.4619, 218.4571, 218.4481, 218.4624, 218.4462, 218.4449, 218.4539, 218.4566, 218.4526, 218.4474, 218.4561, 218.4726, 218.4692, 218.4872, 218.492, 218.4888, 218.4844, 218.4813, 218.486, 218.5089, 218.4445, 218.4864, 218.493, 218.4844, 218.4987, 218.4955, 218.5102, 218.5191, 218.5267, 218.5057, 218.5246, 218.5347, 218.4789, 218.5361, 218.5077, 218.5125, 218.5357, 218.5382, 218.5476, 218.5502, 218.5572, 218.5426, 218.5469, 218.5383, 218.5493, 218.573, 218.5773, 218.5613, 218.5565, 218.5793, 218.5658, 218.5804, 218.5941, 218.5873, 218.5576, 218.5582, 218.5704, 218.5755, 218.5677, 218.6021, 218.5727, 218.5728, 218.5618, 218.5817, 218.5666, 218.603, 218.5891, 218.6073, 218.6098, 218.581, 218.586, 218.6208, 218.587, 218.6085, 218.6313, 218.6373, 218.5942, 205.0363, 31.0056, 11.9238, 12.0028, 11.924, 11.6909, 10.1797, 10.1729, 10.1718, 10.1649, 10.1628, 10.1627, 10.1612, 10.1544, 10.1553, 10.158, 10.1548, 10.167, 10.1604, 10.1619, 10.1521, 10.1493, 10.1405, 10.141, 10.131, 10.1409, 10.1366, 10.1429, 10.1438, 10.1458, 10.1418, 10.1479, 10.148, 10.1467, 10.1425, 10.1489, 10.1535, 10.1568, 10.1538, 10.1569, 10.1547, 10.1544, 10.1579, 10.153, 10.1508, 10.1532, 10.15, 10.1527, 10.1539, 10.1528, 10.1552, 10.151, 10.1547, 10.148, 10.1501, 10.151, 10.15, 10.1486, 10.1506, 10.1514, 10.1501, 10.1504, 10.151, 10.1492, 10.1535, 10.1491, 10.1504, 10.1503, 10.1494, 10.1503, 10.1531, 10.1516, 10.1478, 10.1535, 10.1456, 10.1481, 10.1481, 10.1398, 10.1283, 10.1296, 10.1254, 10.1247, 10.1264, 10.1228, 10.1227, 10.1191, 10.1165, 10.1102, 10.1125, 10.1094, 10.1288, 10.1132, 10.1138, 10.065, 10.0931, 10.085, 10.0943, 10.0942, 10.0926, 10.0939, 10.3468, 10.3016, 10.2969, 10.3118, 10.3176, 10.3223, 10.3207, 10.3234, 10.3232, 10.3275, 10.3274, 10.3333, 10.336, 10.3341, 10.3308, 10.3356, 10.3433, 10.1154, 10.0993, 10.0873, 10.1072, 10.104, 10.1036, 10.1127, 10.1091, 10.1127, 10.1131, 10.1016, 10.1025, 10.1006, 10.1025, 10.1012, 10.1005, 10.1014, 10.1012, 10.1144}
PRES_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
PRES_REL =
  {999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0, 999999.0}
PRES_REL_quality_control =
  {99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99}
DEPTH =
  {206.7933, 206.80286, 206.80956, 206.80609, 206.80609, 206.81602, 206.81271, 206.82242, 206.81575, 206.81256, 206.80286, 206.82257, 206.78978, 206.79631, 206.80623, 206.81602, 206.8094, 206.81602, 206.81602, 206.81595, 206.80623, 206.81602, 206.8129, 206.80968, 206.8129, 206.79976, 206.80286, 206.80319, 206.79973, 206.80968, 206.82242, 206.82593, 206.82257, 206.81929, 206.83566, 206.81595, 206.82582, 206.82565, 206.83237, 206.82912, 206.81602, 206.82912, 206.82912, 206.83247, 206.83585, 206.83247, 206.84206, 206.83533, 206.83557, 206.84221, 206.85175, 206.87488, 206.83885, 206.85513, 206.85187, 206.85498, 206.8454, 206.85513, 206.86478, 206.85513, 206.86478, 206.85513, 206.87785, 206.87466, 206.85513, 206.87466, 206.86145, 206.87778, 206.88458, 206.87466, 206.88791, 206.89761, 206.89095, 206.89095, 206.87785, 206.89761, 206.87785, 206.91722, 206.8943, 206.89095, 206.90736, 206.88765, 206.8943, 206.90388, 206.89413, 206.90065, 206.9009, 206.9009, 206.88765, 206.88763, 206.91385, 206.9009, 206.90729, 206.91057, 206.90404, 206.9204, 206.92679, 206.92377, 206.93333, 206.91075, 206.9301, 206.9301, 206.91695, 206.92679, 206.92024, 206.91695, 206.94337, 206.91695, 206.92024, 206.93333, 206.90729, 206.93028, 206.93341, 206.93996, 206.92995, 206.92024, 206.92995, 206.9266, 206.93988, 206.9266, 206.94319, 206.9431, 206.96597, 206.9431, 206.94641, 206.94641, 206.94975, 206.93968, 206.9365, 206.95277, 206.94958, 206.94608, 206.95932, 206.95277, 206.94948, 206.95596, 206.95932, 206.94958, 206.95944, 206.95296, 206.94958, 206.96571, 206.9692, 206.9824, 206.95627, 206.95932, 206.97586, 206.95612, 206.95944, 206.9596, 206.97234, 206.98538, 206.96251, 206.96284, 206.96579, 206.98538, 206.9853, 206.98207, 206.99178, 206.98877, 206.97891, 206.98538, 206.98538, 206.97552, 206.98877, 206.99544, 207.00514, 206.99211, 206.9853, 206.9853, 207.02142, 206.99196, 206.98538, 206.99524, 206.99193, 207.00179, 207.00514, 206.99847, 207.01479, 207.01158, 206.99193, 206.99847, 206.99524, 206.99832, 206.99832, 206.98877, 207.00491, 207.00491, 207.00818, 207.00491, 207.01479, 206.99178, 206.99516, 206.99496, 207.02795, 207.00163, 207.01794, 207.01813, 207.02464, 207.02464, 207.01828, 207.0146, 207.02448, 207.02464, 207.03769, 207.03432, 207.02795, 207.01488, 207.04405, 207.01488, 207.01479, 207.02127, 207.0278, 207.03113, 207.03102, 207.0443, 207.02795, 207.02127, 207.03102, 207.02467, 207.04086, 207.04405, 207.03432, 207.03102, 207.04094, 207.02762, 207.03432, 207.02115, 207.0474, 207.0375, 207.04405, 207.03087, 207.04405, 207.0439, 207.04086, 207.04094, 207.05394, 207.06686, 207.03766, 207.0439, 207.04094, 207.06049, 207.05394, 207.0735, 207.04405, 207.05045, 207.06049, 207.05707, 207.04721, 207.0603, 207.07, 207.07335, 207.04074, 207.06685, 207.0735, 207.07335, 207.08308, 207.07034, 207.08308, 207.07332, 207.0865, 207.06685, 207.0667, 207.0767, 207.0766, 207.06685, 207.08324, 207.09312, 207.07993, 207.0896, 207.10277, 207.08646, 207.0865, 207.08308, 207.09949, 207.09297, 207.0963, 207.06015, 207.08975, 207.09312, 207.0963, 207.08324, 207.08975, 207.0963, 207.08308, 207.09952, 207.10277, 207.0963, 207.0963, 207.09285, 207.0865, 207.10588, 207.11241, 207.10904, 207.10931, 207.10931, 207.09615, 207.09297, 207.10931, 207.09297, 207.10269, 207.11255, 207.08342, 207.09949, 207.10269, 207.08646, 207.11255, 207.0896, 207.11577, 207.1025, 207.10606, 207.10606, 207.0963, 207.09294, 207.10277, 207.09952, 207.10931, 207.10269, 207.08658, 207.10904, 207.09297, 207.10588, 207.10606, 207.10277, 207.11269, 207.1224, 207.10269, 207.09285, 207.10269, 207.10606, 207.10931, 207.09615, 207.08975, 207.10277, 207.09949, 207.10269, 207.09933, 207.09933, 207.09297, 207.09952, 207.0963, 207.08308, 207.0963, 207.10916, 207.0766, 207.10606, 207.10277, 207.10916, 207.07977, 207.10606, 207.10269, 207.10269, 207.09294, 207.09596, 207.11241, 207.08646, 207.09596, 207.0863, 207.10277, 207.11592, 207.09285, 207.09949, 207.10931, 207.0963, 207.10622, 207.09285, 207.10606, 207.10269, 207.0896, 207.09285, 207.09615, 207.08975, 207.08942, 207.09297, 207.09312, 207.0766, 207.07977, 207.08324, 207.07683, 207.07996, 207.07332, 207.08646, 207.08308, 207.08308, 207.07, 207.07034, 207.07977, 207.06361, 207.07016, 207.0767, 207.0667, 207.07034, 207.08342, 207.06049, 207.0767, 207.07993, 207.05707, 207.06049, 207.07034, 207.06049, 207.04074, 207.0506, 207.04713, 207.06697, 207.04721, 207.04721, 207.05699, 207.04086, 207.0474, 207.05727, 207.0439, 207.03413, 207.0541, 207.04405, 207.04405, 207.0278, 207.04405, 207.03432, 207.0345, 207.03087, 207.03102, 207.02448, 207.0181, 207.04086, 207.03114, 207.03113, 207.02142, 207.00839, 207.02467, 207.00806, 207.01141, 207.01158, 207.01479, 207.01158, 207.00491, 206.99496, 207.00163, 207.00179, 207.01479, 207.00163, 206.98862, 207.00502, 206.99847, 206.99832, 206.99866, 206.99866, 206.9853, 206.97903, 206.99516, 206.98877, 206.98877, 206.98558, 206.96579, 206.9692, 206.9824, 206.9853, 206.96284, 206.96597, 206.97234, 206.96613, 206.96613, 206.96579, 206.97586, 206.96597, 206.95944, 206.95627, 206.95944, 206.95277, 206.95932, 206.9365, 206.94641, 206.94948, 206.94641, 206.92995, 206.94641, 206.93333, 206.93968, 206.9365, 206.93015, 206.9431, 206.9266, 206.94623, 206.9204, 206.93683, 206.92995, 206.93333, 206.92024, 206.9137, 206.92355, 206.91057, 206.90388, 206.91678, 206.90404, 206.91057, 206.89413, 206.89413, 206.9137, 206.8974, 206.90068, 206.90736, 206.87117, 206.9137, 206.8974, 206.90068, 206.89113, 206.8974, 206.89413, 206.88109, 206.89413, 206.89761, 206.89413, 206.87466, 206.89761, 206.87785, 206.88765, 206.8908, 206.87466, 206.85513, 206.87785, 206.87138, 206.8682, 206.86166, 206.89095, 206.87466, 206.86478, 206.86145, 206.8682, 206.86827, 206.86478, 206.85823, 206.85823, 206.85202, 206.86177, 206.84874, 206.8615, 206.84554, 206.86166, 206.85495, 206.85187, 206.85857, 206.85823, 206.86177, 206.85841, 206.83885, 206.83237, 206.85202, 206.84206, 206.84554, 206.84892, 206.83247, 206.83875, 206.83885, 206.83907, 206.82896, 206.84521, 206.83557, 206.82896, 206.83247, 206.82582, 206.83235, 206.81602, 206.83237, 206.81271, 206.81929, 206.82896, 206.80286, 206.81256, 206.82242, 206.82257, 206.80623, 206.82582, 206.79646, 206.8094, 206.8129, 206.81602, 206.7933, 206.78993, 206.79631, 206.79631, 206.79951, 206.78339, 206.79984, 206.80968, 206.78023, 206.79315, 206.78677, 206.81929, 206.76367, 206.77686, 206.79315, 206.78993, 206.77356, 206.79312, 206.76367, 206.78691, 206.79646, 206.78023, 206.78993, 206.79004, 206.78339, 206.78323, 206.77702, 206.78023, 206.77374, 206.7702, 206.78023, 206.77356, 206.76735, 206.75412, 206.76735, 206.76047, 206.76701, 206.74428, 206.75761, 206.74757, 206.75412, 206.77065, 206.75728, 206.76059, 206.76059, 206.74757, 206.74773, 206.75761, 206.76074, 206.75394, 206.74428, 206.7542, 206.74438, 206.74113, 206.75761, 206.74438, 206.75713, 206.75746, 206.75728, 206.74739, 206.73802, 206.7379, 206.73448, 206.75394, 206.74773, 206.74438, 206.73793, 206.73438, 206.75093, 206.75073, 206.75095, 206.74442, 206.75095, 206.74438, 206.7379, 206.73769, 206.74757, 206.74757, 206.73802, 206.74773, 206.74773, 206.73448, 206.7313, 206.7542, 206.75073, 206.7542, 206.74757, 206.74442, 206.73793, 206.74757, 206.74103, 206.74442, 206.73132, 206.7313, 206.73448, 206.76059, 206.74455, 206.76399, 206.74442, 206.76059, 206.75095, 206.73438, 206.74739, 206.76059, 206.75073, 206.76399, 206.77054, 206.76701, 206.75412, 206.76714, 206.75728, 206.76714, 206.76714, 206.77374, 206.76714, 206.77054, 206.77383, 206.76059, 206.75728, 206.77702, 206.76399, 206.77702, 206.76059, 206.78038, 206.7933, 206.77356, 206.78357, 206.76389, 206.7641, 206.76701, 206.75728, 206.76367, 206.77383, 206.76059, 206.77383, 206.76398, 206.75713, 206.77054, 206.76389, 206.77686, 206.76714, 206.76714, 206.77702, 206.76714, 206.77374, 206.78023, 206.78677, 206.76059, 206.77037, 206.78677, 206.7933, 206.78339, 206.76714, 206.79004, 206.7767, 206.78978, 206.7801, 206.78023, 206.79315, 206.79312, 206.79646, 206.79976, 206.78323, 206.77686, 206.79659, 206.80295, 206.8129, 206.79973, 206.79659, 206.79951, 206.78658, 206.80319, 206.79984, 206.80295, 206.81622, 206.80638, 206.8094, 206.80295, 206.80295, 206.81595, 206.83557, 206.80956, 206.81944, 206.82257, 206.80968, 206.81622, 206.80956, 206.82593, 206.80956, 206.82593, 206.8129, 206.81595, 206.81595, 206.82257, 206.81271, 206.80623, 206.80956, 206.83235, 206.82257, 206.82257, 206.82912, 206.83247, 206.82257, 206.8191, 206.83566, 206.85202, 206.8486, 206.8454, 206.83247, 206.82582, 206.84206, 206.8322, 206.83557, 206.83533, 206.86177, 206.83875, 206.83247, 206.84221, 206.83907, 206.85187, 206.84221, 206.83237, 206.84843, 206.83885, 206.83875, 206.85814, 206.8486, 206.84874, 206.84874, 206.85841, 206.86478, 206.86496, 206.86177, 206.8715, 206.86827, 206.87138, 206.87785, 206.86478, 206.86478, 206.87459, 206.87454, 206.88112, 206.8844, 206.87785, 206.8682, 206.87805, 206.8844, 206.88425, 206.86478, 206.8844, 206.8974, 206.88112, 206.88127, 206.8943, 206.90404, 206.88458, 206.89749, 206.89444, 206.89413, 206.90388, 206.88791, 206.88791, 206.90736, 206.90388, 206.90404, 206.90416, 206.90065, 206.90729, 206.90416, 206.8943, 206.9137, 206.9009, 206.91357, 206.90736, 206.90404, 206.91385, 206.89413, 206.91042, 206.93028, 206.9266, 206.91711, 206.91722, 206.92332, 206.94319, 206.93683, 206.94974, 206.92348, 206.93333, 206.92679, 206.93028, 206.93674, 206.94975, 206.94641, 206.93333, 206.95296, 206.92355, 206.9365, 206.93968, 206.95296, 206.95944, 206.94641, 206.93996, 206.94958, 206.95944, 206.93988, 206.9365, 206.94975, 206.9367, 206.96579, 206.95277, 206.95944, 206.96597, 206.96266, 206.96266, 206.96597, 206.96266, 206.97891, 206.95612, 206.96933, 206.97903, 206.95932, 206.97876, 206.97552, 206.99193, 206.99193, 206.9824, 206.97552, 206.98558, 207.00163, 206.98877, 207.00502, 206.98877, 206.99866, 207.00179, 206.99832, 207.01158, 206.98877, 207.00839, 207.00818, 206.99524, 206.99178, 207.00491, 207.00839, 207.00502, 207.01488, 207.01794, 207.00491, 207.02795, 207.00504, 207.00806, 207.00839, 207.01141, 207.02127, 207.00163, 207.00502, 207.01155, 207.00839, 207.00818, 207.01794, 207.04086, 207.02127, 207.01158, 207.01828, 207.03102, 207.01141, 207.02127, 207.04086, 207.03413, 207.0345, 207.0506, 207.02475, 207.03102, 207.0443, 207.01794, 207.03432, 207.03769, 207.04405, 207.0603, 207.03769, 207.05072, 207.0278, 207.04721, 207.03741, 207.04721, 207.0474, 207.04439, 207.0603, 207.0474, 207.0375, 207.05394, 207.0767, 207.08342, 207.05699, 207.05045, 207.0767, 207.06361, 207.08658, 207.0735, 207.0766, 207.08324, 207.07016, 207.05394, 207.0603, 207.0603, 207.06685, 207.0896, 207.08308, 207.07335, 207.08658, 207.08324, 207.07993, 207.0735, 207.08975, 207.0963, 207.08658, 207.08324, 207.08308, 207.0865, 207.09952, 207.10606, 207.11255, 207.09297, 207.10916, 207.10269, 207.08658, 207.09949, 207.08646, 207.11269, 207.10588, 207.10931, 207.11577, 207.11255, 207.0896, 207.10277, 207.11577, 207.11577, 207.1223, 207.11908, 207.10606, 207.10606, 207.10588, 207.1224, 207.10916, 207.11592, 207.11241, 207.10916, 207.10269, 207.10606, 207.10269, 207.12563, 207.12895, 207.11592, 207.10606, 207.12215, 207.11559, 207.12213, 207.12529, 207.11559, 207.1223, 207.12544, 207.1223, 207.1224, 207.1223, 207.13216, 207.1223, 207.1223, 207.1287, 207.13199, 207.1223, 207.13199, 207.1223, 207.12563, 207.13216, 207.12544, 207.13216, 207.11577, 207.15176, 207.13216, 207.11227, 207.13199, 207.1223, 207.12868, 207.13216, 207.12563, 207.10916, 207.13853, 207.11241, 207.14172, 207.13864, 207.1189, 207.11227, 207.13199, 207.10931, 207.13864, 207.11241, 207.1224, 207.12878, 207.10916, 207.11255, 207.10606, 207.10269, 207.11577, 207.11241, 207.11592, 207.12895, 207.12215, 207.11592, 207.1224, 207.11577, 207.10916, 207.11577, 207.12213, 207.10916, 207.11923, 207.11559, 207.12895, 207.10916, 207.10916, 207.10588, 207.10606, 207.11255, 207.09952, 207.11577, 207.1189, 207.09933, 207.0963, 207.09615, 207.1025, 207.10606, 207.09285, 207.10606, 207.09949, 207.1189, 207.09952, 207.11577, 207.1189, 207.1223, 207.08011, 207.08942, 207.0896, 207.10269, 207.09933, 207.10269, 207.08324, 207.07016, 207.10269, 207.07996, 207.07335, 207.07332, 207.08011, 207.07, 207.09285, 207.08011, 207.06049, 207.06361, 207.07996, 207.06361, 207.07034, 207.07332, 207.05376, 207.07335, 207.06697, 207.06697, 207.05394, 207.05072, 207.0766, 207.04755, 207.04405, 207.05394, 207.0443, 207.04721, 207.04721, 207.04721, 207.04086, 207.02795, 207.04721, 207.02448, 207.01794, 207.00818, 207.02127, 207.02464, 207.01479, 207.01479, 206.98862, 207.00502, 206.99193, 207.00514, 206.99193, 206.98862, 207.00179, 206.99847, 206.99211, 206.98222, 206.98877, 206.99178, 206.98889, 206.97903, 206.98207, 206.98538, 206.97574, 206.96251, 206.96933, 206.95932, 206.96579, 206.9596, 206.96266, 206.94958, 206.95612, 206.95627, 206.95296, 206.9364, 206.95296, 206.92995, 206.94656, 206.93333, 206.94974, 206.9367, 206.9365, 206.92024, 206.91042, 206.92679, 206.90404, 206.92024, 206.9204, 206.90388, 206.9137, 206.90404, 206.91406, 206.91075, 206.90388, 206.91711, 206.91711, 206.8974, 206.8844, 206.89749, 206.88765, 206.88425, 206.89761, 206.88112, 206.8844, 206.86804, 206.88127, 206.88127, 206.87138, 206.86496, 206.86478, 206.8484, 206.85841, 206.83885, 206.85187, 206.86827, 206.86478, 206.84193, 206.84554, 206.85529, 206.84874, 206.84221, 206.83237, 206.84892, 206.83885, 206.82884, 206.82565, 206.83585, 206.83247, 206.82896, 206.83557, 206.81944, 206.82582, 206.82896, 206.81944, 206.79646, 206.80623, 206.80621, 206.81622, 206.82257, 206.79312, 206.80621, 206.78023, 206.78658, 206.79984, 206.80286, 206.78323, 206.79631, 206.77037, 206.78658, 206.78993, 206.79004, 206.77054, 206.7865, 206.76714, 206.77037, 206.77356, 206.77374, 206.76399, 206.78023, 206.74757, 206.7801, 206.77686, 206.75412, 206.77374, 206.76735, 206.77054, 206.76735, 206.74739, 206.76735, 206.77374, 206.76389, 206.75073, 206.73448, 206.76399, 206.75743, 206.76059, 206.73448, 206.74428, 206.75093, 206.74773, 206.74442, 206.73122, 206.74773, 206.74773, 206.73463, 206.73448, 206.74438, 206.71812, 206.72467, 206.73448, 206.72478, 206.71173, 206.7214, 206.73476, 206.71812, 206.7184, 206.72156, 206.7085, 206.70181, 206.71487, 206.69537, 206.72156, 206.7085, 206.69211, 206.7281, 206.71829, 206.7053, 206.7053, 206.7085, 206.70518, 206.7085, 206.71173, 206.69856, 206.68912, 206.70518, 206.69565, 206.7085, 206.7087, 206.69884, 206.68884, 206.70518, 206.68245, 206.7087, 206.69884, 206.69211, 206.7087, 206.6859, 206.6792, 206.70181, 206.68245, 206.7053, 206.68893, 206.69229, 206.70552, 206.68893, 206.69229, 206.68893, 206.69884, 206.70518, 206.71504, 206.70518, 206.69864, 206.70203, 206.69856, 206.7087, 206.71191, 206.70181, 206.7053, 206.70181, 206.71504, 206.71828, 206.7281, 206.7214, 206.74739, 206.7313, 206.74757, 206.72467, 206.74113, 206.73802, 206.72795, 206.73463, 206.74757, 206.73448, 206.74442, 206.73122, 206.73448, 206.75412, 206.75412, 206.75412, 206.76399, 206.76389, 206.76059, 206.75412, 206.75073, 206.74773, 206.76399, 206.73769, 206.75412, 206.76399, 206.76399, 206.77383, 206.77065, 206.77037, 206.7542, 206.75728, 206.76367, 206.77374, 206.76398, 206.76047, 206.7641, 206.77054, 206.76059, 206.77702, 206.77065, 206.77054, 206.77374, 206.76735, 206.75728, 206.76399, 206.76398, 206.77374, 206.77686, 206.7767, 206.78023, 206.77686, 206.76389, 206.7801, 206.78339, 206.76714, 206.76714, 206.77065, 206.78691, 206.77686, 206.78323, 206.77356, 206.78993, 206.78357, 206.76701, 206.78677, 206.79004, 206.77383, 206.78993, 206.78677, 206.78323, 206.7933, 206.7866, 206.80319, 206.78357, 206.78993, 206.79315, 206.79315, 206.79659, 206.79984, 206.79659, 206.80968, 206.80286, 206.80319, 206.79984, 206.81602, 206.79303, 206.7933, 206.79315, 206.79303, 206.80621, 206.8094, 206.79984, 206.8094, 206.81929, 206.81944, 206.8094, 206.80956, 206.81944, 206.81929, 206.81622, 206.81602, 206.81595, 206.82565, 206.82242, 206.83235, 206.8223, 206.82896, 206.84554, 206.83907, 206.83566, 206.83907, 206.84554, 206.8258, 206.83907, 206.83557, 206.82242, 206.83533, 206.83557, 206.84206, 206.83885, 206.85187, 206.85175, 206.83533, 206.84206, 206.85187, 206.8486, 206.8486, 206.85823, 206.85823, 206.8486, 206.85513, 206.8486, 206.85841, 206.86177, 206.8682, 206.86827, 206.87466, 206.86496, 206.86827, 206.8682, 206.88127, 206.87778, 206.87138, 206.87785, 206.87785, 206.8715, 206.87805, 206.87778, 206.8682, 206.89095, 206.8844, 206.87466, 206.89095, 206.8682, 206.88776, 206.87778, 206.87785, 206.91075, 206.89761, 206.88127, 206.9009, 206.8943, 206.90068, 206.90736, 206.90388, 206.90068, 206.90416, 206.91057, 206.90404, 206.8908, 206.91075, 206.91385, 206.91057, 206.90703, 206.9009, 206.90703, 206.91711, 206.91695, 206.93333, 206.9137, 206.91357, 206.91711, 206.92377, 206.91357, 206.9367, 206.92694, 206.92679, 206.92355, 206.92348, 206.92694, 206.92679, 206.9365, 206.92332, 206.93321, 206.92995, 206.93321, 206.93968, 206.93988, 206.92995, 206.93321, 206.94623, 206.9431, 206.9266, 206.93988, 206.93968, 206.9431, 206.93321, 206.9364, 206.92679, 206.92355, 206.93321, 206.92355, 206.91695, 206.9137, 206.90388, 206.92355, 206.93015, 206.93321, 206.92024, 206.92995, 206.92995, 206.92995, 206.93321, 206.93028, 206.9365, 206.93321, 206.9431, 206.93968, 206.95277, 206.92995, 206.9266, 206.9365, 206.94623, 206.93683, 206.94974, 206.94641, 206.92679, 206.92995, 206.93321, 206.9431, 206.94958, 206.96281, 206.95296, 206.94656, 206.94641, 206.93341, 206.9364, 206.95612, 206.9431, 206.9432, 206.95944, 206.95612, 206.93321, 206.9432, 206.93988, 206.94958, 206.95296, 206.95277, 206.95296, 206.9692, 206.99193, 206.99524, 206.9853, 206.99193, 207.00163, 206.99178, 207.00163, 207.00839, 206.99832, 207.01158, 207.0181, 206.99832, 207.0181, 207.00818, 207.01158, 207.00151, 207.00502, 207.00163, 206.99496, 207.02127, 207.0181, 207.03769, 207.0146, 207.02448, 207.02115, 207.02762, 207.03413, 207.03114, 207.0443, 207.0474, 207.04094, 207.0375, 207.02762, 207.02795, 207.03741, 207.0443, 207.04094, 207.0345, 207.03784, 207.0474, 207.03413, 207.0345, 207.03413, 207.03769, 207.03114, 207.04405, 207.03769, 207.04755, 207.06032, 207.05394, 207.06346, 207.05394, 207.06685, 207.07332, 207.0638, 207.0735, 207.06361, 207.0767, 207.08342, 207.08646, 207.07996, 207.08342, 207.08324, 207.0896, 207.0963, 207.08975, 207.08975, 207.08975, 207.08975, 207.09312, 207.10916, 207.09615, 207.09933, 207.09952, 207.11255, 207.10916, 207.10606, 207.10606, 207.12213, 207.11592, 207.11559, 207.1223, 207.11241, 207.11577, 207.1223, 207.11577, 207.13864, 207.13515, 207.12868, 207.13533, 207.12868, 207.12868, 207.1223, 207.13853, 207.13533, 207.1485, 207.13853, 207.13853, 207.12868, 207.14516, 207.13184, 207.14516, 207.14497, 207.15813, 207.13853, 207.15143, 207.1679, 207.13834, 207.17451, 207.1615, 207.1646, 207.15813, 207.17769, 207.16785, 207.18423, 207.17758, 207.18413, 207.16452, 207.1615, 207.1876, 207.1876, 207.16478, 207.18744, 207.18423, 207.1876, 207.18423, 207.18744, 207.19061, 207.17433, 207.20044, 207.18727, 207.19398, 207.19731, 207.19382, 207.19061, 207.21368, 207.20699, 207.19731, 207.19077, 207.20699, 207.20384, 207.19731, 207.20384, 207.20355, 207.19716, 207.21353, 207.20699, 207.2068, 207.2068, 207.20032, 207.20699, 207.20699, 207.20714, 207.20714, 207.21368, 207.21341, 207.21341, 207.20044, 207.19716, 207.22008, 207.21672, 207.21341, 207.2068, 207.21693, 207.21353, 207.22333, 207.21341, 207.21341, 207.21693, 207.22318, 207.22008, 207.22643, 207.21353, 207.21672, 207.23314, 207.22008, 207.22661, 207.20714, 207.22643, 207.24298, 207.23631, 207.21341, 207.23314, 207.22643, 207.22008, 207.22661, 207.21024, 207.21008, 207.22987, 207.22333, 207.22015, 207.22333, 207.21988, 207.22633, 207.21988, 207.22318, 207.22318, 207.22333, 207.22995, 207.21024, 207.21988, 207.22342, 207.21024, 207.21988, 207.22676, 207.21024, 207.22342, 207.21024, 207.19382, 207.20062, 207.20032, 207.20699, 207.20044, 207.197, 207.20044, 207.19382, 207.19382, 207.18744, 207.19382, 207.20044, 207.18413, 207.20396, 207.18423, 207.17769, 207.17438, 207.1679, 207.19077, 207.17418, 207.1484, 207.1646, 207.15813, 207.17451, 207.1646, 207.1679, 207.14833, 207.15176, 207.14488, 207.15495, 207.13184, 207.15495, 207.12895, 207.12563, 207.12563, 207.11908, 207.12895, 207.11255, 207.10269, 207.12563, 207.10931, 207.11241, 207.11577, 207.11255, 207.09952, 207.07977, 207.10269, 207.1025, 207.08308, 207.07993, 207.10269, 207.09952, 207.08975, 207.07, 207.08308, 207.08975, 207.08011, 207.07034, 207.08658, 207.0766, 207.07335, 207.07034, 207.06049, 207.06697, 207.05072, 207.05707, 207.05072, 207.02762, 207.0443, 207.02475, 207.02448, 207.01155, 207.00839, 207.02127, 207.00491, 207.00839, 207.01158, 207.00818, 206.9985, 206.99496, 207.01155, 206.98862, 206.98207, 206.98207, 206.97267, 206.9824, 206.99866, 206.97574, 206.97258, 206.97234, 206.96933, 206.95305, 206.95932, 206.95612, 206.9367, 206.95296, 206.94623, 206.9431, 206.94958, 206.93028, 206.92332, 206.92694, 206.92694, 206.9301, 206.92995, 206.92694, 206.93341, 206.90736, 206.8943, 206.90729, 206.9137, 206.90404, 206.89761, 206.9009, 206.89749, 206.88094, 206.87805, 206.88127, 206.8844, 206.8844, 206.86166, 206.87466, 206.87138, 206.8682, 206.8682, 206.86166, 206.8715, 206.85529, 206.85187, 206.83875, 206.8486, 206.83237, 206.83885, 206.82884, 206.82912, 206.82593, 206.8293, 206.82242, 206.82582, 206.83237, 206.82275, 206.82582, 206.80956, 206.8191, 206.80968, 206.79976, 206.7801, 206.81276, 206.79631, 206.80968, 206.80295, 206.79631, 206.79659, 206.78993, 206.76714, 206.80295, 206.78993, 206.76701, 206.77686, 206.7801, 206.77686, 206.77686, 206.77054, 206.77383, 206.76399, 206.76735, 206.76714, 206.76059, 206.76389, 206.76047, 206.75713, 206.76059, 206.76389, 206.74438, 206.75743, 206.75073, 206.7641, 206.74438, 206.74428, 206.75093, 206.74428, 206.73448, 206.72795, 206.73793, 206.73463, 206.73448, 206.73122, 206.73476, 206.72156, 206.7281, 206.74438, 206.72823, 206.73149, 206.72495, 206.7281, 206.7085, 206.70503, 206.72156, 206.70518, 206.7184, 206.72156, 206.7053, 206.69548, 206.71487, 206.71173, 206.69238, 206.70203, 206.69211, 206.71191, 206.70518, 206.70181, 206.69864, 206.6792, 206.69229, 206.69864, 206.70181, 206.6891, 206.68893, 206.68245, 206.70218, 206.68893, 206.67592, 206.69229, 206.68575, 206.67255, 206.68245, 206.66939, 206.68575, 206.68556, 206.68575, 206.69238, 206.68884, 206.68245, 206.68231, 206.68245, 206.68575, 206.67592, 206.68893, 206.68231, 206.69229, 206.68893, 206.67255, 206.68884, 206.68575, 206.68245, 206.70518, 206.6761, 206.6891, 206.68893, 206.69229, 206.68245, 206.67903, 206.67903, 206.70203, 206.69211, 206.69211, 206.69864, 206.69229, 206.70218, 206.69566, 206.68575, 206.69229, 206.69211, 206.71191, 206.69891, 206.70842, 206.7053, 206.71504, 206.71487, 206.70203, 206.71173, 206.70181, 206.7085, 206.70203, 206.71173, 206.70203, 206.72156, 206.7053, 206.71191, 206.71828, 206.71828, 206.70552, 206.69548, 206.71158, 206.73149, 206.71828, 206.7214, 206.7214, 206.72174, 206.71487, 206.73463, 206.72156, 206.72475, 206.71828, 206.72795, 206.72795, 206.73463, 206.73448, 206.7281, 206.7281, 206.72156, 206.74739, 206.73793, 206.73122, 206.74103, 206.73476, 206.7379, 206.74103, 206.73802, 206.74086, 206.7379, 206.74103, 206.75746, 206.7313, 206.73802, 206.74442, 206.73122, 206.77065, 206.75093, 206.73793, 206.75394, 206.74739, 206.76735, 206.75412, 206.75095, 206.74739, 206.76389, 206.76735, 206.77037, 206.75746, 206.77037, 206.77686, 206.77702, 206.77037, 206.7801, 206.78677, 206.77356, 206.78658, 206.7767, 206.77702, 206.77702, 206.79646, 206.78339, 206.79659, 206.78023, 206.78677, 206.7933, 206.7933, 206.78677, 206.79646, 206.78993, 206.79646, 206.78978, 206.79984, 206.80295, 206.78677, 206.80638, 206.80623, 206.79312, 206.79984, 206.80286, 206.81944, 206.82275, 206.81595, 206.80638, 206.81276, 206.81929, 206.80956, 206.81276, 206.81602, 206.81944, 206.82242, 206.83566, 206.8258, 206.83907, 206.82896, 206.85529, 206.83557, 206.83882, 206.83907, 206.86177, 206.8486, 206.84874, 206.85202, 206.85187, 206.85841, 206.84874, 206.86166, 206.85513, 206.86166, 206.8454, 206.85823, 206.86478, 206.8682, 206.86166, 206.87117, 206.86469, 206.88127, 206.88127, 206.86478, 206.87117, 206.87805, 206.89761, 206.88765, 206.89113, 206.88776, 206.89749, 206.89113, 206.9009, 206.88765, 206.89095, 206.90753, 206.90068, 206.89413, 206.90404, 206.90416, 206.90068, 206.90404, 206.90729, 206.9137, 206.92024, 206.90388, 206.90416, 206.91711, 206.92006, 206.91057, 206.9137, 206.91695, 206.92355, 206.9137, 206.92355, 206.92006, 206.93996, 206.9301, 206.91678, 206.9301, 206.91711, 206.92006, 206.9266, 206.9301, 206.9301, 206.9301, 206.93988, 206.9301, 206.91357, 206.93333, 206.92694, 206.9301, 206.9367, 206.92377, 206.93028, 206.9301, 206.94974, 206.9365, 206.93988, 206.94623, 206.94319, 206.94319, 206.95277, 206.94958, 206.96597, 206.94975, 206.96266, 206.94623, 206.95932, 206.95296, 206.96579, 206.96579, 206.94948, 206.9693, 206.95596, 206.96912, 206.94958, 206.95627, 206.94641, 206.96266, 206.96579, 206.9692, 206.96597, 206.95612, 206.97574, 206.95917, 206.9824, 206.97903, 206.98862, 206.98877, 206.97585, 206.98222, 206.97922, 206.9692, 206.97234, 206.98207, 206.99211, 206.97903, 206.98222, 206.98877, 206.98207, 206.98558, 206.98538, 206.97891, 206.99866, 206.99524, 206.98877, 206.98862, 207.00179, 206.99524, 207.00818, 207.01167, 206.98862, 206.99544, 206.99178, 206.99832, 207.01155, 207.01479, 207.01158, 207.02464, 207.02467, 206.99847, 207.01479, 207.00806, 207.00818, 207.00491, 207.00818, 206.99516, 207.02464, 207.01479, 207.0278, 207.0146, 207.02448, 207.04086, 207.02464, 207.04074, 207.02795, 207.03769, 207.04086, 207.02467, 207.04086, 207.03113, 207.0375, 207.05072, 207.03113, 207.0603, 207.04405, 207.03087, 207.04405, 207.0439, 207.05072, 207.05707, 207.06049, 207.06685, 207.05072, 207.0603, 207.0603, 207.06685, 207.06685, 207.08308, 207.08658, 207.0767, 207.0766, 207.09642, 207.0963, 207.0865, 207.0865, 207.08293, 207.09952, 207.11592, 207.10277, 207.10269, 207.11241, 207.09952, 207.1224, 207.12563, 207.13216, 207.1189, 207.1223, 207.11908, 207.12895, 207.12544, 207.11577, 207.12213, 207.11577, 207.13199, 207.13199, 207.15176, 207.1484, 207.13853, 207.13853, 207.14516, 207.13515, 207.13853, 207.14516, 207.14516, 207.14833, 207.15495, 207.15495, 207.15813, 207.15797, 207.1646, 207.16785, 207.18085, 207.17758, 207.17451, 207.17769, 207.1615, 207.19095, 207.17451, 207.19398, 207.17769, 207.18413, 207.19061, 207.19716, 207.19716, 207.18085, 207.19409, 207.19077, 207.20699, 207.19077, 207.20062, 207.19731, 207.19716, 207.19382, 207.20699, 207.21033, 207.22015, 207.21024, 207.22342, 207.22643, 207.22318, 207.22661, 207.21988, 207.21988, 207.23297, 207.24937, 207.24268, 207.2362, 207.22987, 207.24268, 207.23969, 207.25253, 207.2362, 207.24283, 207.25253, 207.25278, 207.26227, 207.25926, 207.25572, 207.2556, 207.26881, 207.25587, 207.2787, 207.26552, 207.26897, 207.26552, 207.26552, 207.28171, 207.27855, 207.27216, 207.27888, 207.2849, 207.29176, 207.2948, 207.2919, 207.29497, 207.2915, 207.29814, 207.2948, 207.30466, 207.31436, 207.30151, 207.308, 207.30135, 207.30135, 207.2916, 207.30788, 207.2948, 207.3045, 207.29832, 207.32108, 207.31427, 207.30135, 207.29802, 207.32419, 207.32095, 207.31436, 207.32419, 207.31755, 207.31137, 207.3146, 207.3177, 207.31436, 207.32419, 207.32108, 207.33058, 207.32747, 207.3308, 207.33401, 207.32419, 207.32762, 207.32762, 207.31755, 207.31783, 207.32735, 207.32108, 207.33092, 207.30788, 207.32108, 207.308, 207.3177, 207.30151, 207.33733, 207.32443, 207.3178, 207.3339, 207.31427, 207.32443, 207.30481, 207.308, 207.30788, 207.31136, 207.32095, 207.30162, 207.30481, 207.3177, 207.30788, 207.2819, 207.31783, 207.30466, 207.308, 207.2915, 207.28838, 207.29176, 207.30162, 207.27873, 207.29497, 207.28523, 207.26227, 207.27216, 207.26881, 207.26572, 207.27206, 207.26227, 207.27216, 207.25587, 207.26567, 207.25572, 207.25926, 207.25587, 207.25587, 207.24606, 207.24617, 207.24283, 207.25572, 207.23936, 207.23952, 207.25572, 207.2365, 207.23297, 207.22987, 207.2362, 207.24268, 207.23631, 207.2068, 207.23631, 207.22643, 207.21988, 207.21341, 207.19061, 207.19716, 207.21368, 207.20044, 207.197, 207.18744, 207.18413, 207.18106, 207.18106, 207.19409, 207.1679, 207.18727, 207.16785, 207.17467, 207.1646, 207.16132, 207.15813, 207.14813, 207.13853, 207.13853, 207.13518, 207.1417, 207.12868, 207.13199, 207.13864, 207.12578, 207.13216, 207.12544, 207.11923, 207.11908, 207.11592, 207.10916, 207.10931, 207.09615, 207.10588, 207.09952, 207.08011, 207.08342, 207.07977, 207.0766, 207.07683, 207.0735, 207.0667, 207.05699, 207.08011, 207.06361, 207.0506, 207.04713, 207.05045, 207.04405, 207.04094, 207.02448, 207.02464, 207.02115, 207.01479, 207.01155, 207.02142, 207.00179, 207.01488, 207.00839, 206.99193, 206.99832, 206.97234, 206.97574, 206.97891, 206.97891, 206.97891, 206.9692, 206.96266, 206.95944, 206.96579, 206.9693, 206.93996, 206.95296, 206.95277, 206.94656, 206.93321, 206.92355, 206.9367, 206.93028, 206.93683, 206.92355, 206.92355, 206.91695, 206.91711, 206.90416, 206.90729, 206.90703, 206.90404, 206.8943, 206.90065, 206.8943, 206.88127, 206.87466, 206.88127, 206.8844, 206.86145, 206.87785, 206.86166, 206.88763, 206.86478, 206.86166, 206.86478, 206.86478, 206.84521, 206.83885, 206.83875, 206.85187, 206.84892, 206.82912, 206.82912, 206.82884, 206.81926, 206.79976, 206.80638, 206.81622, 206.80638, 206.78339, 206.81271, 206.81276, 206.80319, 206.82582, 206.80621, 206.78677, 206.79004, 206.78339, 206.77686, 206.7866, 206.77702, 206.78357, 206.75394, 206.78023, 206.77054, 206.76399, 206.75728, 206.74428, 206.75761, 206.74103, 206.76047, 206.74103, 206.73793, 206.75093, 206.7641, 206.7641, 206.72467, 206.72795, 206.74438, 206.70842, 206.74455, 206.71828, 206.71191, 206.71173, 206.71173, 206.7214, 206.73448, 206.71828, 206.7379, 206.7281, 206.70203, 206.72174, 206.70842, 206.7085, 206.69864, 206.70203, 206.69864, 206.7085, 206.69211, 206.68245, 206.69884, 206.69884, 206.70181, 206.68893, 206.69864, 206.6792, 206.67903, 206.68575, 206.68245, 206.66618, 206.6761, 206.68884, 206.69864, 206.69565, 206.66939, 206.66628, 206.66946, 206.68245, 206.65308, 206.67265, 206.66628, 206.66618, 206.67265, 206.6466, 206.69229, 206.66284, 206.66628, 206.67265, 206.66628, 206.66312, 206.6563, 206.66922, 206.65645, 206.64642, 206.64339, 206.6563, 206.65976, 206.66284, 206.6563, 206.6563, 206.65321, 206.6594, 206.65321, 206.65009, 206.65648, 206.65321, 206.65645, 206.65657, 206.65614, 206.66628, 206.6563, 206.66312, 206.67577, 206.6466, 206.65308, 206.67592, 206.66284, 206.67265, 206.68575, 206.68231, 206.6695, 206.6594, 206.66284, 206.6695, 206.68259, 206.69864, 206.6792, 206.67265, 206.68884, 206.69238, 206.68245, 206.66594, 206.68256, 206.69566, 206.69548, 206.68556, 206.69229, 206.68575, 206.69238, 206.68575, 206.69211, 206.69864, 206.7085, 206.69856, 206.70518, 206.69196, 206.71523, 206.70181, 206.71173, 206.7087, 206.70842, 206.73448, 206.71504, 206.72495, 206.7085, 206.72495, 206.72495, 206.7184, 206.7379, 206.71173, 206.72156, 206.73769, 206.74739, 206.72467, 206.73122, 206.74113, 206.72467, 206.74113, 206.7511, 206.74428, 206.7542, 206.74739, 206.73448, 206.73793, 206.76398, 206.73793, 206.75728, 206.75743, 206.74757, 206.75095, 206.75394, 206.75394, 206.76735, 206.77383, 206.76059, 206.78357, 206.77037, 206.77702, 206.78357, 206.77686, 206.75095, 206.80319, 206.78357, 206.77356, 206.79976, 206.80638, 206.8129, 206.79659, 206.82896, 206.8094, 206.79312, 206.79631, 206.80609, 206.79951, 206.8094, 206.83237, 206.81271, 206.8191, 206.83566, 206.8191, 206.8322, 206.81929, 206.82896, 206.83557, 206.8191, 206.8129, 206.83566, 206.8486, 206.83907, 206.84874, 206.85529, 206.8486, 206.82582, 206.8486, 206.85187, 206.82896, 206.87805, 206.8615, 206.85175, 206.86166, 206.87459, 206.8844, 206.87785, 206.86496, 206.8715, 206.88127, 206.87459, 206.88458, 206.85175, 206.86496, 206.87138, 206.87466, 206.88776, 206.85495, 206.8974, 206.88136, 206.87488, 206.88763, 206.89761, 206.89413, 206.91406, 206.90736, 206.8844, 206.88776, 206.9009, 206.8908, 206.92006, 206.90404, 206.90404, 206.90729, 206.90729, 206.90388, 206.93333, 206.9301, 206.93341, 206.9137, 206.90068, 206.8974, 206.92995, 206.92024, 206.90736, 206.93996, 206.9266, 206.89749, 206.90388, 206.91695, 206.92355, 206.9266, 206.91711, 206.9137, 206.9367, 206.94975, 206.9431, 206.93683, 206.93996, 206.93321, 206.95932, 206.93341, 206.92679, 206.92024, 206.94319, 206.95932, 206.97574, 206.96579, 206.96266, 206.94958, 206.9431, 206.95296, 206.9596, 206.9563, 206.96912, 206.96933, 206.94623, 206.9596, 206.93968, 206.92348, 206.92348, 206.9365, 206.94974, 206.95612, 206.94974, 206.95944, 206.95944, 206.95296, 206.98207, 206.98222, 206.93968, 206.96579, 206.97221, 206.97552, 206.98538, 206.9985, 206.9692, 206.97891, 206.96912, 206.99193, 206.97903, 206.97922, 206.95262, 206.98222, 206.97876, 206.96912, 206.97891, 206.96912, 206.97891, 207.00179, 206.97876, 207.00514, 206.99196, 207.00491, 206.99211, 206.99178, 206.9853, 206.99178, 206.98207, 206.99524, 206.98222, 206.99211, 207.00502, 206.99516, 207.00179, 206.98877, 207.01813, 207.00514, 207.00818, 207.01813, 206.99524, 207.01488, 207.02448, 207.01828, 207.00491, 207.02475, 207.00851, 206.99832, 206.99832, 206.99496, 207.00504, 207.02464, 207.01813, 207.00806, 207.01158, 207.01813, 207.01158, 206.98843, 207.0278, 207.01488, 207.00163, 207.0443, 207.01479, 207.01479, 207.03769, 207.03741, 207.00839, 207.0181, 207.02762, 207.05376, 207.02434, 207.0375, 207.02762, 207.0146, 207.02115, 207.03432, 207.04074, 207.03741, 207.03102, 207.04074, 207.05394, 207.06697, 207.03741, 207.0474, 207.03741, 207.06685, 207.0375, 207.0375, 207.0541, 207.05394, 207.05394, 207.07977, 207.0767, 207.06685, 207.06712, 207.07332, 207.07977, 207.08658, 207.09285, 207.08942, 207.10277, 207.10606, 207.0896, 207.11255, 207.09615, 207.0896, 207.10269, 207.1025, 207.11592, 207.11908, 207.12563, 207.11592, 207.1224, 207.12878, 207.13518, 207.13853, 207.13199, 207.1417, 207.14516, 207.12878, 207.13533, 207.16132, 207.14488, 207.14186, 207.14497, 207.15477, 207.14828, 207.16165, 207.17769, 207.1548, 207.15825, 207.15825, 207.1646, 207.17451, 207.18423, 207.18413, 207.19398, 207.20044, 207.17467, 207.17438, 207.20396, 207.19382, 207.1876, 207.19398, 207.20044, 207.2068, 207.19716, 207.21672, 207.22015, 207.21024, 207.21696, 207.22661, 207.21988, 207.22972, 207.22972, 207.23314, 207.22008, 207.24927, 207.23969, 207.22318, 207.24937, 207.25253, 207.23297, 207.23952, 207.24617, 207.24954, 207.24606, 207.26227, 207.25253, 207.25572, 207.2459, 207.2626, 207.26552, 207.27191, 207.26215, 207.28198, 207.27206, 207.27206, 207.28198, 207.28838, 207.29178, 207.29814, 207.28838, 207.29507, 207.30466, 207.30481, 207.28838, 207.30151, 207.2916, 207.31116, 207.28171, 207.31116, 207.31116, 207.31137, 207.30788, 207.32095, 207.32419, 207.32074, 207.32095, 207.32744, 207.3177, 207.33401, 207.31116, 207.35359, 207.33058, 207.34056, 207.33058, 207.34381, 207.34381, 207.33746, 207.34372, 207.34071, 207.34056, 207.36006, 207.34705, 207.3308, 207.33719, 207.3569, 207.36664, 207.35008, 207.36009, 207.36983, 207.3666, 207.35342, 207.37311, 207.3569, 207.36644, 207.35342, 207.36009, 207.36644, 207.37619, 207.36676, 207.36664, 207.35342, 207.37619, 207.36328, 207.36664, 207.36644, 207.3829, 207.39615, 207.37965, 207.37637, 207.38602, 207.36345, 207.3991, 207.3666, 207.37619, 207.39594, 207.36664, 207.38927, 207.38945, 207.37326, 207.37651, 207.36983, 207.3731, 207.38945, 207.36983, 207.39275, 207.36964, 207.37938, 207.37299, 207.38945, 207.37651, 207.37938, 207.3731, 207.36676, 207.37651, 207.36328, 207.38626, 207.37965, 207.36998, 207.36998, 207.3666, 207.36983, 207.33733, 207.3536, 207.3568, 207.36009, 207.36009, 207.33058, 207.35042, 207.3308, 207.35359, 207.33058, 207.34705, 207.34071, 207.32735, 207.3308, 207.32762, 207.32744, 207.33719, 207.31108, 207.3045, 207.31137, 207.33401, 207.2915, 207.2948, 207.3045, 207.2916, 207.30135, 207.31137, 207.308, 207.308, 207.28171, 207.29176, 207.28528, 207.2919, 207.27518, 207.26572, 207.26863, 207.27855, 207.24927, 207.25244, 207.26242, 207.26881, 207.24617, 207.2658, 207.24283, 207.22643, 207.22643, 207.23282, 207.22972, 207.21341, 207.23314, 207.22015, 207.2362, 207.21672, 207.21368, 207.19052, 207.2068, 207.18423, 207.22015, 207.20062, 207.17758, 207.21353, 207.18413, 207.18423, 207.17114, 207.1679, 207.15477, 207.15813, 207.1615, 207.17451, 207.16132, 207.15143, 207.1548, 207.13853, 207.13834, 207.1485, 207.10277, 207.14186, 207.10588, 207.12563, 207.09933, 207.10916, 207.11577, 207.10916, 207.10277, 207.09615, 207.09615, 207.06686, 207.09297, 207.0766, 207.07332, 207.07683, 207.07016, 207.06346, 207.06032, 207.05394, 207.05727, 207.02448, 207.02762, 207.03769, 207.03102, 207.03114, 207.02127, 207.0278, 207.01479, 206.99832, 207.01479, 207.01794, 206.99832, 206.98538, 207.00151, 206.99866, 206.95944, 206.99832, 206.98207, 206.97234, 206.96266, 206.98222, 206.95296, 206.95296, 206.97221, 206.95612, 206.9596, 206.94623, 206.93333, 206.9365, 206.9431, 206.93321, 206.93333, 206.9301, 206.91695, 206.9204, 206.91385, 206.90404, 206.90388, 206.91711, 206.88425, 206.89113, 206.87466, 206.8844, 206.88748, 206.86478, 206.87488, 206.87466, 206.88127, 206.85823, 206.85823, 206.8486, 206.83885, 206.86166, 206.83585, 206.85187, 206.8486, 206.83557, 206.84521, 206.82565, 206.82896, 206.80956, 206.81929, 206.78993, 206.82257, 206.8191, 206.7865, 206.77383, 206.80286, 206.78978, 206.7702, 206.77383, 206.77686, 206.76714, 206.77054, 206.78023, 206.77702, 206.75412, 206.75412, 206.75095, 206.73438, 206.75073, 206.7511, 206.73438, 206.74103, 206.75761, 206.74442, 206.71487, 206.73448, 206.71504, 206.74113, 206.72495, 206.71812, 206.7281, 206.71504, 206.69548, 206.71504, 206.71828, 206.69884, 206.69548, 206.71487, 206.69864, 206.7087, 206.68575, 206.70181, 206.69884, 206.69229, 206.67903, 206.6859, 206.6859, 206.68245, 206.68245, 206.67265, 206.69238, 206.71176, 206.67903, 206.66594, 206.68259, 206.68893, 206.68556, 206.6596, 206.6761, 206.67607, 206.66939, 206.69884, 206.66939, 206.67935, 206.69229, 206.66284, 206.66293, 206.68556, 206.68884, 206.68912, 206.6594, 206.67592, 206.68256, 206.67935, 206.68245, 206.6594, 206.67282, 206.6594, 206.6859, 206.67903, 206.67265, 206.67255, 206.67265, 206.65308, 206.68575, 206.66284, 206.66594, 206.66594, 206.67265, 206.6792, 206.6594, 206.64995, 206.66939, 206.6594, 206.66618, 206.66618, 206.67282, 206.67935, 206.68575, 206.6792, 206.6792, 206.6695, 206.65308, 206.68245, 206.66312, 206.65308, 206.6762, 206.66284, 206.6792, 206.66939, 206.67255, 206.66618, 206.67255, 206.68245, 206.66628, 206.68556, 206.68256, 206.68556, 206.68245, 206.68575, 206.69238, 206.67592, 206.69211, 206.69891, 206.69884, 206.70203, 206.69864, 206.68912, 206.69229, 206.70181, 206.69884, 206.71504, 206.69211, 206.7053, 206.7053, 206.69548, 206.7085, 206.71812, 206.71828, 206.72495, 206.71504, 206.71828, 206.71812, 206.73463, 206.71828, 206.73149, 206.74442, 206.73463, 206.73463, 206.7379, 206.72795, 206.74438, 206.74455, 206.7214, 206.74438, 206.74757, 206.74113, 206.74757, 206.73793, 206.74428, 206.75073, 206.76059, 206.76047, 206.75728, 206.76399, 206.76735, 206.77374, 206.75073, 206.75728, 206.76399, 206.75095, 206.78339, 206.75412, 206.76389, 206.75412, 206.78677, 206.78691, 206.7933, 206.79315, 206.7933, 206.80319, 206.79312, 206.80638, 206.78339, 206.80621, 206.82242, 206.82257, 206.82257, 206.82896, 206.82593, 206.81595, 206.81602, 206.82582, 206.81256, 206.82912, 206.83557, 206.84521, 206.83885, 206.84206, 206.8486, 206.84221, 206.8322, 206.83557, 206.83237, 206.84221, 206.83875, 206.85841, 206.86469, 206.8454, 206.8682, 206.86496, 206.85823, 206.86827, 206.86166, 206.86177, 206.87778, 206.87488, 206.87138, 206.87778, 206.8908, 206.88425, 206.87805, 206.8715, 206.87785, 206.88127, 206.8715, 206.8844, 206.87138, 206.86827, 206.90404, 206.88109, 206.89113, 206.8908, 206.89761, 206.89113, 206.89095, 206.8974, 206.90068, 206.90404, 206.8974, 206.89761, 206.91711, 206.91385, 206.90736, 206.91695, 206.89761, 206.90736, 206.92694, 206.91695, 206.92694, 206.91711, 206.91075, 206.9137, 206.92377, 206.9266, 206.93683, 206.92006, 206.91695, 206.9301, 206.93015, 206.92355, 206.9137, 206.92679, 206.90068, 206.9204, 206.91357, 206.91042, 206.92006, 206.93988, 206.9365, 206.93341, 206.9431, 206.93988, 206.93333, 206.94337, 206.92679, 206.93988, 206.95627, 206.95944, 206.94641, 206.94641, 206.95944, 206.93988, 206.93988, 206.94974, 206.9364, 206.95612, 206.94623, 206.9367, 206.94293, 206.94319, 206.92995, 206.94623, 206.93968, 206.95612, 206.94623, 206.94641, 206.93341, 206.9365, 206.93968, 206.94958, 206.95296, 206.92694, 206.9365, 206.94958, 206.94948, 206.94293, 206.95296, 206.93028, 206.93988, 206.9364, 206.91711, 206.9364, 206.93968, 206.94975, 206.95596, 206.9596, 206.95612, 206.95627, 206.95612, 206.93341, 206.9365, 206.94958, 206.94641, 206.96266, 206.9563, 206.95932, 206.95627, 206.95612, 206.95612, 206.95596, 206.95612, 206.95917, 206.94958, 206.96571, 206.97234, 206.94623, 206.94641, 206.94641, 206.95627, 206.95612, 206.9853, 206.98538, 206.97876, 206.9596, 206.97574, 206.98222, 206.95305, 206.96912, 206.96266, 206.96266, 206.9692, 206.97876, 206.99544, 207.00502, 206.9853, 206.98877, 206.98207, 206.99193, 206.98222, 207.00504, 206.99832, 206.99524, 206.99866, 206.99847, 206.99524, 207.02127, 207.02475, 207.00491, 207.00514, 207.0146, 207.00491, 207.01813, 207.02464, 207.03087, 207.02142, 207.01479, 207.02142, 207.02467, 207.0345, 207.02464, 207.02127, 207.03113, 207.04405, 207.05394, 207.04755, 207.02115, 207.05376, 207.04755, 207.0443, 207.0443, 207.05379, 207.0474, 207.06049, 207.0603, 207.0638, 207.05394, 207.05394, 207.06049, 207.0735, 207.09615, 207.06361, 207.07016, 207.07034, 207.05707, 207.06361, 207.0735, 207.0667, 207.0667, 207.0735, 207.0896, 207.0896, 207.1025, 207.07332, 207.08658, 207.0896, 207.1189, 207.10606, 207.10916, 207.11923, 207.1223, 207.10904, 207.10588, 207.11908, 207.1417, 207.14186, 207.13199, 207.13548, 207.14516, 207.15813, 207.13853, 207.14828, 207.1484, 207.15176, 207.15158, 207.17114, 207.17418, 207.16452, 207.15813, 207.15797, 207.18085, 207.18423, 207.17769, 207.18727, 207.19398, 207.20369, 207.18396, 207.19382, 207.19409, 207.19382, 207.21988, 207.20369, 207.21024, 207.21353, 207.21341, 207.22015, 207.21353, 207.22995, 207.21693, 207.22643, 207.25253, 207.243, 207.25278, 207.23952, 207.25926, 207.23936, 207.25587, 207.25253, 207.27206, 207.28516, 207.25253, 207.2459, 207.24283, 207.25587, 207.26242, 207.25899, 207.2787, 207.25899, 207.25572, 207.27206, 207.26863, 207.28838, 207.27206, 207.2916, 207.31137, 207.3178, 207.29814, 207.29802, 207.29178, 207.30466, 207.29497, 207.31116, 207.32108, 207.308, 207.31783, 207.32771, 207.3177, 207.32095, 207.30481, 207.32735, 207.3308, 207.31783, 207.3341, 207.31436, 207.33733, 207.33733, 207.32443, 207.34726, 207.3502, 207.33719, 207.34381, 207.33719, 207.34726, 207.36345, 207.36009, 207.36317, 207.35042, 207.3339, 207.34705, 207.36676, 207.35994, 207.36644, 207.36328, 207.36964, 207.39275, 207.38278, 207.37637, 207.37965, 207.34705, 207.38602, 207.38626, 207.38945, 207.35657, 207.38306, 207.3666, 207.37953, 207.37311, 207.37965, 207.37619, 207.39902, 207.39615, 207.3603, 207.37637, 207.40262, 207.3829, 207.3829, 207.39902, 207.38626, 207.37938, 207.38278, 207.38626, 207.38278, 207.39275, 207.37962, 207.37651, 207.37637, 207.37283, 207.37283, 207.37651, 207.39275, 207.37637, 207.38945, 207.37962, 207.4025, 207.36983, 207.38306, 207.3991, 207.38602, 207.37637, 207.38602, 207.39594, 207.37965, 207.37326, 207.36328, 207.36964, 207.36009, 207.36998, 207.38945, 207.37965, 207.36006, 207.34038, 207.35657, 207.3568, 207.35994, 207.36328, 207.34706, 207.3568, 207.35342, 207.36345, 207.3537, 207.3536, 207.34053, 207.35042, 207.35008, 207.33398, 207.3241, 207.34053, 207.33058, 207.32443, 207.3341, 207.3341, 207.31436, 207.33058, 207.308, 207.32419, 207.31116, 207.32095, 207.30788, 207.3241, 207.32744, 207.30466, 207.31137, 207.2983, 207.2948, 207.29802, 207.2916, 207.26897, 207.2948, 207.26881, 207.2948, 207.27216, 207.2819, 207.2556, 207.27206, 207.24937, 207.24927, 207.25899, 207.24617, 207.21988, 207.2362, 207.24617, 207.23631, 207.22333, 207.21024, 207.22995, 207.22342, 207.22333, 207.20699, 207.21353, 207.20384, 207.21024, 207.19398, 207.18434, 207.17418, 207.20699, 207.18744, 207.15825, 207.18423, 207.16478, 207.17099, 207.1679, 207.14201, 207.15176, 207.1484, 207.13533, 207.13216, 207.14186, 207.12563, 207.11559, 207.12578, 207.10916, 207.12544, 207.1025, 207.08324, 207.09967, 207.09285, 207.0863, 207.0865, 207.09312, 207.07996, 207.08342, 207.04074, 207.06346, 207.05394, 207.0474, 207.05045, 207.03413, 207.04086, 207.02762, 207.02127, 207.00491, 207.01794, 207.00502, 206.99866, 207.02434, 207.02795, 206.99211, 206.99196, 206.98558, 206.98538, 206.97267, 206.9692, 206.97574, 206.97574, 206.98889, 206.95612, 206.95612, 206.94623, 206.9204, 206.94623, 206.9365, 206.91057, 206.9367, 206.9236, 206.9367, 206.89749, 206.90404, 206.9204, 206.90404, 206.9009, 206.88748, 206.90068, 206.90736, 206.90416, 206.87785, 206.88425, 206.89113, 206.86511, 206.86478, 206.85187, 206.85187, 206.83885, 206.86478, 206.85187, 206.85187, 206.81929, 206.83875, 206.80623, 206.83885, 206.81595, 206.81602, 206.82593, 206.83585, 206.82565, 206.78993, 206.81622, 206.78993, 206.78978, 206.79346, 206.7865, 206.76714, 206.78339, 206.77037, 206.79315, 206.77054, 206.78357, 206.76701, 206.7801, 206.76059, 206.76047, 206.75746, 206.75073, 206.73793, 206.75073, 206.74757, 206.73149, 206.7511, 206.69864, 206.72495, 206.70181, 206.73149, 206.70842, 206.71829, 206.69211, 206.71487, 206.71158, 206.7053, 206.69548, 206.70181, 206.69856, 206.6792, 206.69211, 206.7053, 206.68575, 206.71504, 206.6859, 206.68893, 206.6792, 206.67592, 206.68245, 206.68245, 206.6695, 206.67592, 206.68245, 206.67265, 206.66618, 206.6594, 206.65645, 206.68575, 206.6761, 206.66284, 206.66972, 206.67265, 206.69238, 206.66939, 206.67265, 206.63353, 206.66284, 206.65645, 206.66296, 206.66628, 206.6466, 206.64975, 206.67265, 206.63675, 206.65657, 206.63675, 206.6399, 206.63014, 206.65308, 206.65645, 206.63684, 206.63362, 206.64006, 206.63362, 206.6399, 206.62067, 206.63048, 206.65009, 206.61722, 206.63335, 206.67265, 206.6303, 206.61722, 206.63362, 206.6466, 206.61722, 206.6236, 206.6303, 206.6466, 206.66284, 206.65009, 206.64034, 206.65308, 206.6596, 206.65009, 206.65648, 206.6399, 206.63675, 206.65321, 206.6467, 206.6563, 206.63362, 206.6466, 206.64323, 206.64034, 206.6792, 206.65645, 206.65614, 206.66618, 206.63675, 206.66312, 206.6594, 206.6695, 206.67282, 206.65321, 206.6499, 206.67282, 206.67265, 206.67592, 206.6859, 206.67577, 206.67903, 206.69211, 206.68259, 206.6859, 206.6761, 206.69238, 206.69211, 206.70503, 206.69884, 206.68893, 206.67607, 206.70842, 206.71191, 206.73132, 206.70181, 206.69884, 206.71523, 206.7053, 206.71158, 206.7085, 206.7053, 206.71173, 206.73463, 206.73448, 206.71828, 206.69548, 206.7085, 206.72495, 206.73463, 206.72122, 206.7313, 206.7281, 206.73476, 206.73448, 206.75073, 206.73448, 206.73448, 206.72795, 206.74428, 206.77686, 206.77374, 206.76735, 206.78023, 206.76399, 206.76059, 206.77383, 206.77374, 206.77054, 206.76735, 206.77374, 206.78658, 206.78677, 206.80295, 206.80956, 206.80638, 206.79976, 206.79984, 206.80295, 206.8293, 206.76059, 206.80295, 206.80956, 206.79976, 206.81602, 206.8094, 206.82582, 206.8322, 206.84206, 206.82257, 206.84221, 206.85187, 206.79312, 206.8484, 206.82242, 206.82565, 206.85187, 206.85175, 206.86496, 206.86478, 206.87138, 206.85495, 206.85814, 206.85175, 206.86827, 206.89113, 206.8943, 206.87459, 206.87138, 206.89761, 206.87778, 206.89413, 206.91057, 206.90753, 206.87813, 206.87466, 206.88776, 206.89095, 206.88112, 206.9204, 206.89113, 206.89113, 206.88136, 206.89749, 206.88458, 206.9204, 206.90056, 206.92355, 206.92348, 206.90099, 206.90068, 206.93321, 206.90068, 206.92694, 206.94293, 206.95296, 206.91057, 193.45847, 20.724241, 1.7790508, 1.8580271, 1.7755916, 1.5455393, 0.048100777, 0.041229334, 0.037779845, 0.030908957, 0.030922484, 0.030923048, 0.027475799, 0.020604327, 0.024054931, 0.02749548, 0.020602083, 0.034352846, 0.02748027, 0.030927526, 0.020618968, 0.017178984, 0.01032045, 0.010317653, -0.0034481469, 0.010318215, 0.0034309581, 0.010305252, 0.010300217, 0.013744684, 0.0068557486, 0.013731166, 0.013730604, 0.017195303, 0.013764919, 0.020638647, 0.024066793, 0.024046533, 0.020607684, 0.020588549, 0.020602643, 0.020604327, 0.027496042, 0.017156504, 0.013713161, 0.024068473, 0.017175065, 0.017158184, 0.020607123, 0.017157625, 0.02751292, 0.020625122, 0.020602643, 0.013730604, 0.017174508, 0.020625122, 0.017175065, 0.013727247, 0.013714277, 0.020622887, 0.017174508, 0.017172825, 0.020625122, 0.017179541, 0.024066793, 0.0171801, 0.017172825, 0.017173385, 0.017178422, 0.017173385, 0.02406903, 0.020621765, 0.013731718, 0.024066793, 0.013745801, 0.013730043, 0.013730043, 0.0034112828, -0.0068878243, -0.0034385535, -0.010326383, -0.010322465, -0.006875435, -0.010310078, -0.010309517, -0.013744162, -0.017184408, -0.024058748, -0.024073372, -0.024054268, -0.00343408, -0.02062074, -0.017167551, -0.068716735, -0.034322266, -0.048099674, -0.037787262, -0.037786704, -0.037776023, -0.041241575, 0.21298085, 0.16486904, 0.16144165, 0.17863238, 0.18550919, 0.18893662, 0.18549, 0.185473, 0.1889316, 0.1923612, 0.19236177, 0.19923793, 0.19922097, 0.19923344, 0.19925387, 0.20268065, 0.21300237, -0.020634802, -0.03090389, -0.04811428, -0.024040215, -0.02747712, -0.03093142, -0.020617943, -0.027509153, -0.020617943, -0.02062018, -0.030918486, -0.02746698, -0.034369446, -0.02746698, -0.03091625, -0.034368884, -0.030917373, -0.03091625, -0.017170908}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
}
