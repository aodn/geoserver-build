netcdf file-45.nc {
  dimensions:
    DEPTH = 48;
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852, 22572.18258101852}
TEMP =
  {19.5733, 19.5656, 19.5607, 19.5141, 19.4961, 19.471, 19.4423, 19.4242, 19.4195, 19.4134, 19.4043, 19.3981, 19.3931, 19.3849, 19.3813, 19.3796, 19.3783, 19.3763, 19.3746, 19.3737, 19.3731, 19.3721, 19.3694, 19.3687, 19.3682, 19.3667, 19.3662, 19.3659, 19.3657, 19.3658, 19.3658, 19.3658, 19.3652, 19.3646, 19.3629, 19.3581, 19.3558, 19.3529, 19.3485, 19.3317, 19.2854, 19.2625, 19.2393, 19.2164, 19.2073, 19.2039, 19.2015, 19.2015}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
