netcdf file-44.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (47 currently)
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705, 22545.094953703705}
TEMP =
  {20.0698, 20.0698, 20.0571, 20.0529, 20.0454, 20.0365, 20.0314, 20.025, 20.0239, 20.024, 20.0221, 20.0219, 20.0224, 20.0228, 20.0231, 20.0239, 20.0232, 20.0228, 20.021, 20.0198, 20.0185, 20.017, 20.015, 20.0126, 20.0096, 20.0065, 20.0055, 20.0051, 20.0057, 20.0041, 20.0031, 20.0034, 20.0038, 20.0042, 20.0043, 20.0045, 20.0046, 20.0047, 20.0047, 20.0049, 20.005, 20.0048, 20.0049, 20.0052, 20.0059, 20.0081, 99999.0}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
