netcdf file-84.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334, 23178.480208333334}
TEMP =
  {27.0166, 27.046, 27.0455, 27.0451, 27.0479, 27.0474, 27.044, 27.0433, 27.0426, 27.0417, 27.0416, 27.0423, 27.0448, 27.0448, 27.0423, 27.0407, 27.0331, 27.0398, 27.0351, 27.0265, 27.0227}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.963, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872}
}
