netcdf file-150.nc {
  dimensions:
    DEPTH = 12;
  variables:
    float LATITUDE(DEPTH=12);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=12);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=12);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=12);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=12);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=12);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184, 21933.049872685184}
TEMP =
  {28.4921, 28.49, 28.4896, 28.4878, 28.4848, 28.4833, 28.483, 28.483, 28.4829, 28.483, 28.4831, 28.4832}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {13.915, 14.909, 15.903, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.854, 24.847}
}
