netcdf file-117.nc {
  dimensions:
    DEPTH = 20;
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037, 22987.93818287037}
TEMP =
  {31.8598, 31.8605, 31.8619, 31.8628, 31.8635, 31.8605, 31.8603, 31.8614, 31.8616, 31.8607, 31.8589, 31.8579, 31.8575, 31.858, 31.8581, 31.8588, 31.8587, 31.8586, 31.8589, 31.8591}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879}
}
