netcdf file-157.nc {
  dimensions:
    DEPTH = 27;
  variables:
    float LATITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=27);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=27);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=27);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=27);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222, 22297.06440972222}
TEMP =
  {29.5591, 29.2427, 29.0595, 29.0059, 29.0366, 29.0655, 29.0812, 29.0893, 29.0985, 29.0892, 29.009, 28.89, 28.7973, 28.7248, 28.6663, 28.639, 28.6243, 28.6184, 28.616, 28.6142, 28.6125, 28.6111, 28.6108, 28.6114, 28.6136, 28.6127, 28.6136}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.957, 7.952, 8.945, 9.94, 10.933, 11.927, 12.921, 13.915, 14.909, 15.902, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835}
}
