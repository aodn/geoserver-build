netcdf file-122.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (21 currently)
  variables:
    float LATITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=21);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=21);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=21);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=21);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556, 22988.123368055556}
TEMP =
  {32.172, 32.1718, 32.1332, 32.0537, 32.0021, 31.9834, 31.9767, 31.9727, 31.9678, 31.9574, 31.9523, 31.9354, 31.9209, 31.911, 31.9022, 31.8977, 31.8955, 31.8939, 31.893, 31.8917, 31.8904}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.965, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.914, 15.908, 16.902, 17.896, 18.891, 19.884, 20.879, 21.873}
}
