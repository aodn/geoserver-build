netcdf file-119.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (20 currently)
  variables:
    float LATITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=20);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=20);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=20);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=20);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625, 22988.0240625}
TEMP =
  {31.9752, 31.9713, 31.9737, 31.9712, 31.9562, 31.9382, 31.9255, 31.9165, 31.9075, 31.8997, 31.8936, 31.8912, 31.8882, 31.885, 31.8776, 31.8739, 31.8742, 31.8725, 31.87, 31.8677}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.989, 2.983, 3.977, 4.971, 5.966, 6.96, 7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.919, 14.913, 15.908, 16.902, 17.896, 18.89, 19.884, 20.879}
}
