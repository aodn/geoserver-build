netcdf file-167.nc {
  dimensions:
    DEPTH = 28;
  variables:
    float LATITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=28);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=28);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=28);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=28);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365, -19.30365}
LONGITUDE =
  {147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391, 147.6391}
TIME =
  {22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964, 22626.127650462964}
TEMP =
  {28.8216, 28.6863, 28.615, 28.571, 28.5316, 28.4942, 28.4296, 28.2762, 28.047, 27.8454, 27.7188, 27.6648, 27.6455, 27.6341, 27.6274, 27.6188, 27.6091, 27.6052, 27.6025, 27.6006, 27.5991, 27.5959, 27.5937, 27.5918, 27.5882, 27.5857, 27.5851, 27.5855}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {0.994, 1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.952, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.903, 16.897, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86, 23.853, 24.847, 25.841, 26.835, 27.829}
}
