netcdf file-49.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (47 currently)
  variables:
    float LATITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=47);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=47);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=47);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=47);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778, 22788.20184027778}
TEMP =
  {22.6215, 22.6269, 22.6274, 22.6272, 22.6267, 22.6247, 22.6128, 22.5881, 22.5483, 22.5183, 22.5021, 22.4919, 22.4839, 22.4692, 22.4497, 22.4313, 22.4212, 22.4125, 22.3957, 22.3857, 22.375, 22.3725, 22.3718, 22.369, 22.3649, 22.3511, 22.3397, 22.339, 22.3368, 22.3351, 22.3336, 22.3339, 22.3334, 22.3305, 22.3295, 22.3295, 22.3292, 22.3291, 22.3285, 22.3277, 22.3272, 22.3264, 22.3266, 22.3268, 22.3268, 22.3271, 22.3275}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
