netcdf file-97.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (13 currently)
  variables:
    float LATITUDE(DEPTH=13);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=13);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=13);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=13);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=13);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=13);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372, -12.3372}
LONGITUDE =
  {130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974, 130.6974}
TIME =
  {22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778, 22658.81402777778}
TEMP =
  {31.5303, 31.5303, 31.534, 31.5394, 31.5403, 31.5414, 31.5416, 31.5416, 31.5416, 31.5403, 31.5391, 31.5378, 31.5365}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {7.954, 8.948, 9.942, 10.937, 11.931, 12.925, 13.92, 14.914, 15.908, 16.902, 17.896, 18.89, 19.885}
}
