netcdf file-158.nc {
  dimensions:
    DEPTH = UNLIMITED;   // (22 currently)
  variables:
    float LATITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=22);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=22);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=22);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=22);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467, -19.303467}
LONGITUDE =
  {147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079, 147.62079}
TIME =
  {22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926, 22327.07550925926}
TEMP =
  {28.7228, 28.715, 28.6996, 28.6692, 28.6359, 28.609, 28.5902, 28.5766, 28.5649, 28.5575, 28.5535, 28.5513, 28.5504, 28.5488, 28.5445, 28.5407, 28.5401, 28.5404, 28.5405, 28.5401, 28.54, 28.5402}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {1.988, 2.982, 3.976, 4.97, 5.964, 6.958, 7.951, 8.945, 9.939, 10.933, 11.927, 12.921, 13.915, 14.909, 15.902, 16.896, 17.89, 18.884, 19.878, 20.872, 21.866, 22.86}
}
