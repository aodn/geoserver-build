netcdf file-15.nc {
  dimensions:
    DEPTH = 43;
  variables:
    float LATITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=43);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=43);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=43);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=43);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93, -33.93}
LONGITUDE =
  {121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85, 121.85}
TIME =
  {22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258, 22808.082071759258}
TEMP =
  {18.1767, 18.1761, 18.1774, 18.1753, 18.1745, 18.1764, 18.1763, 18.1772, 18.1767, 18.1757, 18.1766, 18.1746, 18.1718, 18.1692, 18.1691, 18.1692, 18.1692, 18.169, 18.1691, 18.17, 18.1698, 18.1698, 18.17, 18.1707, 18.1709, 18.1709, 18.1708, 18.1705, 18.17, 18.1711, 18.1706, 18.1708, 18.1712, 18.1716, 18.1727, 18.1728, 18.172, 18.1714, 18.1717, 18.1723, 18.173, 18.173, 18.1716}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0}
}
