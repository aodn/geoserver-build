netcdf file-41.nc {
  dimensions:
    DEPTH = 44;
  variables:
    float LATITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=44);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=44);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=44);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=44);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148, 22452.09741898148}
TEMP =
  {21.2944, 21.3009, 21.3038, 21.3052, 21.3071, 21.3058, 21.3093, 21.3097, 21.3082, 21.2789, 21.2076, 21.1616, 21.1179, 21.0818, 21.0626, 21.0548, 21.046, 21.028, 20.9563, 20.8538, 20.8133, 20.7927, 20.7669, 20.6967, 20.6204, 20.5673, 20.4942, 20.4016, 20.3111, 20.2109, 20.1036, 19.9894, 19.9053, 19.824, 19.7006, 19.6523, 19.6391, 19.6358, 19.6337, 19.6298, 19.627, 19.6241, 19.6237, 19.624}
DEPTH_quality_control =
  {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
DEPTH =
  {4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0}
}
