netcdf file-34.nc {
  dimensions:
    DEPTH = 48;
  variables:
    float LATITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    float LONGITUDE(DEPTH=48);
      :_FillValue = 99999.0f; // float

    double TIME(DEPTH=48);
      :_FillValue = 99999.0; // double
      :units = "days since 1950-01-01 00:00:00 UTC";

    float TEMP(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :example = "examplevalue";

    byte DEPTH_quality_control(DEPTH=48);
      :_FillValue = 0B; // byte

    float DEPTH(DEPTH=48);
      :_FillValue = 99999.0f; // float
      :units = "days since 1950-01-01 00:00:00 UTC";

 data:
LATITUDE =
  {-32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0, -32.0}
LONGITUDE =
  {115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4, 115.4}
TIME =
  {22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223, 22181.199097222223}
TEMP =
  {20.8373, 20.1181, 19.948, 19.9061, 19.8837, 19.8666, 19.8522, 19.8393, 19.8234, 19.8141, 19.8102, 19.8089, 19.805, 19.8008, 19.7935, 19.784, 19.7777, 19.7744, 19.7706, 19.7671, 19.7635, 19.7569, 19.751, 19.7405, 19.7254, 19.7137, 19.7062, 19.7016, 19.7011, 19.7006, 19.6934, 19.6446, 19.5199, 19.2616, 18.9113, 18.6434, 18.4893, 18.2877, 18.1354, 18.0834, 18.0515, 18.0193, 18.0084, 17.9961, 17.9934, 17.9878, 17.9822, 17.9813}
DEPTH_quality_control =
  {4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4}
DEPTH =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0}
}
